#Note:
#IP Version:v0p1
#DK Version:v0p1
SITE  uhd50_CoreSite
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	0.480 BY 3.36 ;
END  uhd50_CoreSite

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AD1V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AD1V1_7TV50 0 0 ;
  SIZE 14.88 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.13 1.91 4.815 2.1 ;
        RECT 4.4 1.91 4.815 2.28 ;
        RECT 6.135 1.41 10.745 1.6 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.84 1.8 7.1 2.32 ;
        RECT 6.84 1.8 9.745 1.99 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 0.32 4.2 1.32 ;
        RECT 0.68 1.13 4.2 1.32 ;
        RECT 3.96 0.32 7.865 0.51 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.525 0.595 12.715 2.43 ;
        RECT 12.525 2 12.84 2.43 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.28 0.56 14.47 2.475 ;
        RECT 14.28 0.56 14.76 0.88 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.595 2.735 1.875 3.48 ;
        RECT 3.355 2.395 3.635 3.48 ;
        RECT 8.12 2.59 8.4 3.48 ;
        RECT 10 2.97 10.28 3.48 ;
        RECT 13.43 2.28 13.665 3.48 ;
        RECT 0 3.24 14.88 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.56 -0.12 1.84 0.93 ;
        RECT 3.315 -0.12 3.595 0.93 ;
        RECT 8.17 -0.12 8.45 0.82 ;
        RECT 10.03 -0.12 10.31 0.43 ;
        RECT 13.38 -0.12 13.66 0.705 ;
        RECT 0 -0.12 14.88 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.205 -0.24 8.735 1.56 ;
        RECT 5.445 -0.24 8.735 1.575 ;
        RECT -0.12 -0.24 15 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.205 3.94 ;
        RECT -0.58 1.56 5.445 3.94 ;
        RECT 8.74 1.46 15.46 3.94 ;
        RECT -0.58 1.575 15.46 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.345 2.785 2.535 ;
      RECT 9.09 2.58 11.19 2.77 ;
      RECT 9.07 0.63 11.275 0.82 ;
      RECT 5.015 0.74 5.295 0.93 ;
      RECT 0.2 1.52 5.245 1.71 ;
      RECT 11.33 1.99 11.52 2.38 ;
      RECT 7.335 2.19 11.52 2.38 ;
      RECT 0.2 0.595 0.39 2.58 ;
      RECT 5.055 0.74 5.245 2.945 ;
      RECT 7.335 2.19 7.525 2.945 ;
      RECT 5.055 2.755 7.525 2.945 ;
      RECT 11.935 0.585 12.125 1.21 ;
      RECT 5.655 1.02 12.125 1.21 ;
      RECT 13.04 1.805 14.04 1.995 ;
      RECT 5.655 0.71 5.845 2.555 ;
      RECT 5.655 2.365 5.935 2.555 ;
      RECT 11.805 1.02 11.995 2.82 ;
      RECT 13.04 1.805 13.23 2.82 ;
      RECT 11.805 2.63 13.23 2.82 ;
  END
END AD1V1_7TV50

MACRO AD1V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AD1V2_7TV50 0 0 ;
  SIZE 16.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.56 2.32 1.8 ;
        RECT 2 1.61 4.755 1.8 ;
        RECT 6.355 1.41 11.06 1.6 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.32 1.8 7.6 2.32 ;
        RECT 7.32 1.8 10.09 1.99 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.68 1.36 ;
        RECT 4.49 0.32 4.68 1.36 ;
        RECT 0.68 1.17 4.68 1.36 ;
        RECT 4.49 0.32 5.915 0.51 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.59 0.64 13.78 2.43 ;
        RECT 13.545 2 13.825 2.43 ;
        RECT 13.59 0.64 13.875 0.83 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 15.29 0.595 15.48 2.475 ;
        RECT 15.29 0.595 15.76 0.84 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.595 2.78 1.875 3.48 ;
        RECT 3.295 2.47 3.575 3.48 ;
        RECT 8.585 2.71 8.865 3.48 ;
        RECT 10.345 2.97 10.625 3.48 ;
        RECT 12.695 2.745 12.93 3.48 ;
        RECT 14.44 2.275 14.675 3.48 ;
        RECT 16.095 2.275 16.375 3.48 ;
        RECT 0 3.24 16.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.645 -0.12 1.925 0.58 ;
        RECT 1.645 -0.12 3.725 0.125 ;
        RECT 3.445 -0.12 3.725 0.815 ;
        RECT 8.385 -0.12 8.665 0.775 ;
        RECT 10.245 -0.12 10.525 0.39 ;
        RECT 12.695 -0.12 12.975 0.75 ;
        RECT 14.495 -0.12 14.775 0.75 ;
        RECT 16.295 -0.12 16.575 0.75 ;
        RECT 0 -0.12 16.8 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.03 -0.24 8.935 1.53 ;
        RECT 5.575 -0.24 8.935 1.575 ;
        RECT -0.12 -0.24 16.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.03 3.94 ;
        RECT -0.58 1.53 5.575 3.94 ;
        RECT 8.935 1.46 17.38 3.94 ;
        RECT -0.58 1.575 17.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.39 2.725 2.58 ;
      RECT 1.1 0.595 1.29 0.97 ;
      RECT 2.59 0.595 2.78 0.97 ;
      RECT 1.1 0.78 2.78 0.97 ;
      RECT 9.285 0.59 11.485 0.78 ;
      RECT 9.435 2.58 11.535 2.77 ;
      RECT 4.995 0.71 5.48 0.9 ;
      RECT 0.2 2 5.185 2.19 ;
      RECT 11.675 1.775 11.865 2.38 ;
      RECT 7.8 2.19 11.865 2.38 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 4.995 0.71 5.185 2.965 ;
      RECT 7.8 2.19 7.99 2.965 ;
      RECT 4.995 2.775 7.99 2.965 ;
      RECT 5.875 1.02 12.34 1.21 ;
      RECT 14.025 1.805 15.05 1.995 ;
      RECT 12.15 0.595 12.34 2.49 ;
      RECT 5.875 0.71 6.065 2.575 ;
      RECT 12.15 2.3 13.345 2.49 ;
      RECT 5.875 2.385 6.405 2.575 ;
      RECT 13.155 2.3 13.345 2.82 ;
      RECT 14.025 1.805 14.215 2.82 ;
      RECT 13.155 2.63 14.215 2.82 ;
  END
END AD1V2_7TV50

MACRO ADH1V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADH1V1_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 0.56 2.76 1.22 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.05 1.85 4.68 2.04 ;
        RECT 4.44 1.85 4.68 2.32 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.335 0.595 0.9 0.84 ;
        RECT 0.71 0.595 0.9 2.475 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.68 0.6 6.87 2.48 ;
        RECT 6.68 0.6 7.255 0.84 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.515 2.675 1.795 3.48 ;
        RECT 3.275 2.33 3.555 3.48 ;
        RECT 5.785 2.28 6.065 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.235 -0.12 1.515 0.765 ;
        RECT 6.12 -0.12 6.355 0.75 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 3.655 -0.24 5.805 1.47 ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.385 3.94 ;
        RECT 5.535 1.46 8.26 3.94 ;
        RECT -0.58 1.47 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.98 0.505 3.17 1.65 ;
      RECT 1.66 1.46 5.53 1.65 ;
      RECT 1.14 1.805 1.85 1.995 ;
      RECT 1.66 1.46 1.85 2.475 ;
      RECT 1.66 2.285 2.705 2.475 ;
      RECT 4.32 0.65 5.92 0.84 ;
      RECT 5.73 0.65 5.92 2.045 ;
      RECT 6.205 1.765 6.395 2.045 ;
      RECT 4.92 1.855 6.395 2.045 ;
      RECT 4.92 1.855 5.11 2.52 ;
  END
END ADH1V1_7TV50

MACRO ADH1V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADH1V2_7TV50 0 0 ;
  SIZE 9.6 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 0.56 3.72 1.26 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.98 1.85 5.64 2.04 ;
        RECT 5.375 1.85 5.64 2.32 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.355 0.6 1.89 0.84 ;
        RECT 1.7 0.6 1.89 2.48 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.11 0.6 8.3 2.48 ;
        RECT 8.11 0.6 8.56 0.84 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.805 2.28 1.085 3.48 ;
        RECT 2.505 2.69 2.785 3.48 ;
        RECT 4.205 2.3 4.485 3.48 ;
        RECT 6.935 2.75 7.215 3.48 ;
        RECT 8.915 2.28 9.195 3.48 ;
        RECT 0 3.24 9.6 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.455 -0.12 0.735 0.765 ;
        RECT 2.255 -0.12 2.535 0.7 ;
        RECT 7.41 -0.12 7.645 0.79 ;
        RECT 9.165 -0.12 9.445 0.735 ;
        RECT 0 -0.12 9.6 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.9 -0.24 5.79 1.53 ;
        RECT -0.12 -0.24 9.72 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.1 3.94 ;
        RECT 6.99 1.46 10.18 3.94 ;
        RECT -0.58 1.53 10.18 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 4.59 0.595 4.78 1.05 ;
      RECT 6.405 0.71 6.685 0.9 ;
      RECT 4.59 0.86 6.595 1.05 ;
      RECT 4 0.545 4.19 1.65 ;
      RECT 6.525 1.37 6.715 1.65 ;
      RECT 2.59 1.46 6.715 1.65 ;
      RECT 2.13 1.81 2.78 2 ;
      RECT 2.59 1.46 2.78 2.475 ;
      RECT 2.59 2.285 3.635 2.475 ;
      RECT 5.535 0.32 7.195 0.51 ;
      RECT 5.445 0.47 5.725 0.66 ;
      RECT 7.005 1.81 7.87 2 ;
      RECT 7.005 0.32 7.195 2.285 ;
      RECT 5.85 2.095 7.195 2.285 ;
      RECT 5.85 2.095 6.04 2.81 ;
  END
END ADH1V2_7TV50

MACRO AND2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.985 1.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.695 1.485 2.28 1.84 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.375 2.23 0.655 3.48 ;
        RECT 1.97 2.885 2.25 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.025 -0.12 2.305 0.835 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.97 0.56 3.16 2.475 ;
        RECT 2.97 0.56 3.24 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.325 0.64 1.46 0.83 ;
      RECT 1.27 1.075 2.68 1.265 ;
      RECT 1.27 0.64 1.46 2.475 ;
  END
END AND2V1_7TV50

MACRO AND2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.18 1.56 3.76 1.81 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.08 2.51 1.365 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.28 0.435 3.48 ;
        RECT 1.855 2.28 2.135 3.48 ;
        RECT 3.555 2.27 3.835 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.72 ;
        RECT 1.955 -0.12 2.235 0.695 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.05 0.56 1.24 2.475 ;
        RECT 1.05 0.56 1.32 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.75 0.64 3.935 0.83 ;
      RECT 1.48 1.805 2.94 1.995 ;
      RECT 2.75 0.64 2.94 2.475 ;
  END
END AND2V2_7TV50

MACRO AND2V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2V4_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.08 1.675 1.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.375 1.8 ;
        RECT 0.745 1.61 3.375 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.27 2.35 0.55 3.48 ;
        RECT 1.97 2.52 2.25 3.48 ;
        RECT 3.67 2.52 3.95 3.48 ;
        RECT 5.37 2.355 5.65 3.48 ;
        RECT 7.07 2.285 7.35 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.22 -0.12 0.5 0.75 ;
        RECT 3.62 -0.12 3.9 0.75 ;
        RECT 5.42 -0.12 5.7 0.625 ;
        RECT 7.22 -0.12 7.5 0.73 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.565 0.595 4.755 1.015 ;
        RECT 4.565 1.965 4.755 2.475 ;
        RECT 5.465 0.825 5.655 2.155 ;
        RECT 4.565 1.965 6.455 2.155 ;
        RECT 6.265 1.965 6.455 2.475 ;
        RECT 6.36 0.56 6.6 1.015 ;
        RECT 4.565 0.825 6.6 1.015 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.965 0.595 2.155 1.22 ;
      RECT 1.965 1.03 3.765 1.22 ;
      RECT 3.575 1.395 4.975 1.585 ;
      RECT 3.575 1.03 3.765 2.32 ;
      RECT 1.165 2.13 3.765 2.32 ;
      RECT 1.165 2.13 1.355 2.48 ;
      RECT 2.865 2.13 3.055 2.48 ;
  END
END AND2V4_7TV50

MACRO AND3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.705 1.075 1.36 1.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.42 1.56 2.02 1.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.335 1.04 2.785 1.36 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.03 2.4 1.31 3.48 ;
        RECT 2.73 2.4 3.01 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.68 -0.12 2.96 0.84 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 0.595 3.815 0.84 ;
        RECT 3.625 0.595 3.815 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.15 1.76 3.34 2.2 ;
      RECT 0.225 2.01 3.34 2.2 ;
      RECT 0.225 0.595 0.415 2.475 ;
      RECT 1.925 2.01 2.115 2.48 ;
  END
END AND3V1_7TV50

MACRO AND3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3V2_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.87 1.04 1.32 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.865 1.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.34 1.04 2.76 1.385 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.695 1.485 3.48 ;
        RECT 2.905 2.695 3.185 3.48 ;
        RECT 4.605 2.28 4.885 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.855 -0.12 3.135 0.705 ;
        RECT 4.655 -0.12 4.935 0.725 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8 0.56 3.99 2.475 ;
        RECT 3.8 0.56 4.2 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.4 0.595 0.59 2.475 ;
      RECT 3.325 1.76 3.515 2.475 ;
      RECT 0.4 2.285 3.515 2.475 ;
  END
END AND3V2_7TV50

MACRO AND3V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3V4_7TV50 0 0 ;
  SIZE 10.56 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.06 1.045 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.06 2.92 1.39 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.695 1.56 5.295 1.8 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.24 2.495 1.52 3.48 ;
        RECT 2.94 2.685 3.22 3.48 ;
        RECT 4.64 2.685 4.92 3.48 ;
        RECT 6.34 2.685 6.62 3.48 ;
        RECT 8.04 2.675 8.32 3.48 ;
        RECT 9.74 2.295 10.02 3.48 ;
        RECT 0 3.24 10.56 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.64 -0.12 4.92 0.76 ;
        RECT 6.44 -0.12 6.72 0.815 ;
        RECT 8.24 -0.12 8.52 0.58 ;
        RECT 10.04 -0.12 10.32 0.745 ;
        RECT 0 -0.12 10.56 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.385 0.595 7.575 0.97 ;
        RECT 8.98 0.78 9.17 2.435 ;
        RECT 7.19 2.235 9.17 2.435 ;
        RECT 9.185 0.56 9.48 0.97 ;
        RECT 7.385 0.78 9.48 0.97 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.965 -0.24 4.715 1.585 ;
        RECT -0.12 -0.24 10.68 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.965 3.94 ;
        RECT 4.715 1.46 11.14 3.94 ;
        RECT -0.58 1.585 11.14 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.435 0.375 4.24 0.565 ;
      RECT 4.05 0.375 4.24 0.955 ;
      RECT 0.435 0.375 0.625 0.86 ;
      RECT 2.295 0.375 2.485 0.86 ;
      RECT 4.05 0.765 4.33 0.955 ;
      RECT 3.15 0.765 3.43 0.955 ;
      RECT 3.24 0.765 3.43 1.345 ;
      RECT 5.585 0.595 5.775 1.345 ;
      RECT 3.24 1.155 5.775 1.345 ;
      RECT 1.35 0.765 1.63 0.955 ;
      RECT 1.44 0.765 1.63 1.995 ;
      RECT 1.44 1.805 2.325 1.995 ;
      RECT 5.535 1.805 7.845 1.995 ;
      RECT 2.135 2.295 5.725 2.485 ;
      RECT 2.135 1.805 2.325 2.6 ;
      RECT 3.835 2.295 4.025 2.6 ;
      RECT 5.535 1.805 5.725 2.6 ;
  END
END AND3V4_7TV50

MACRO AND4V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.52 0.84 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.03 1.86 1.455 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.33 1.49 2.8 1.8 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.945 1.04 3.46 1.32 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.275 0.435 3.48 ;
        RECT 1.855 2.4 2.135 3.48 ;
        RECT 3.615 2.4 3.895 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.495 -0.12 3.775 0.835 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 0.56 4.7 0.88 ;
        RECT 4.51 0.56 4.7 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.195 0.64 1.24 0.83 ;
      RECT 4.035 1.76 4.225 2.2 ;
      RECT 1.05 2.01 4.225 2.2 ;
      RECT 1.05 0.64 1.24 2.475 ;
      RECT 2.75 2.01 2.94 2.475 ;
  END
END AND4V1_7TV50

MACRO AND4V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4V2_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.52 0.84 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.075 1.84 1.525 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 1.56 2.8 1.8 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 0.94 3.34 1.32 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.245 0.435 3.48 ;
        RECT 1.855 2.68 2.135 3.48 ;
        RECT 3.555 2.68 3.835 3.48 ;
        RECT 5.255 2.28 5.535 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.505 -0.12 3.785 0.745 ;
        RECT 5.305 -0.12 5.585 0.715 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.45 0.56 4.64 2.475 ;
        RECT 4.44 0.56 4.68 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.205 0.64 1.24 0.83 ;
      RECT 1.05 0.64 1.24 2.475 ;
      RECT 3.975 1.76 4.165 2.475 ;
      RECT 1.05 2.285 4.165 2.475 ;
  END
END AND4V2_7TV50

MACRO AO112V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO112V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.48 1.52 0.93 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.72 1.8 2.32 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.125 1.76 3.315 2.32 ;
        RECT 3 2 3.315 2.32 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.475 1.56 2.8 2.005 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.615 2.23 3.895 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.885 -0.12 2.165 0.83 ;
        RECT 1.885 -0.12 3.965 0.125 ;
        RECT 3.685 -0.12 3.965 0.83 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.51 0.6 4.7 2.475 ;
        RECT 4.4 0.6 4.865 0.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.28 2.28 0.47 2.865 ;
      RECT 2 2.285 2.19 2.865 ;
      RECT 0.28 2.675 2.19 2.865 ;
      RECT 0.185 0.64 1.32 0.83 ;
      RECT 2.83 0.595 3.02 1.31 ;
      RECT 4.105 1.03 4.295 1.31 ;
      RECT 1.13 1.12 4.295 1.31 ;
      RECT 1.13 0.64 1.32 2.475 ;
  END
END AO112V1_7TV50

MACRO AO112V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO112V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 1.04 0.89 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 2.01 1.84 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.16 1.56 3.76 1.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.46 1.76 2.65 2.28 ;
        RECT 2.46 1.975 2.8 2.28 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.54 2.265 3.82 3.48 ;
        RECT 5.24 2.285 5.52 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.89 -0.12 2.17 0.715 ;
        RECT 3.69 -0.12 3.97 0.715 ;
        RECT 1.89 -0.12 5.77 0.125 ;
        RECT 5.49 -0.12 5.77 0.725 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.635 0.595 4.825 2.76 ;
        RECT 4.39 2.52 4.825 2.76 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.24 2.75 2.22 2.94 ;
      RECT 0.19 0.64 1.325 0.83 ;
      RECT 2.835 0.595 3.025 1.265 ;
      RECT 1.135 1.075 4.345 1.265 ;
      RECT 1.135 0.64 1.325 2.475 ;
  END
END AO112V2_7TV50

MACRO AO12V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO12V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.515 1.52 1.8 2.04 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.84 1.63 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.31 1.52 2.76 1.995 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.78 2.355 3.06 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.23 -0.12 0.51 0.83 ;
        RECT 2.83 -0.12 3.11 0.875 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.675 0.56 3.865 2.475 ;
        RECT 3.675 0.56 4.2 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.275 2.355 0.465 3.025 ;
      RECT 1.975 2.355 2.165 3.025 ;
      RECT 0.275 2.835 2.165 3.025 ;
      RECT 1.975 0.595 2.165 1.31 ;
      RECT 3.25 1.03 3.44 1.31 ;
      RECT 1.125 1.12 3.44 1.31 ;
      RECT 1.125 1.12 1.315 2.475 ;
  END
END AO12V1_7TV50

MACRO AO12V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO12V2_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.695 1.56 2.32 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.995 1.405 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 1.72 2.76 2.32 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.965 2.26 3.2 3.48 ;
        RECT 4.62 2.26 4.9 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.37 -0.12 0.65 0.765 ;
        RECT 2.97 -0.12 3.25 0.765 ;
        RECT 4.77 -0.12 5.05 0.73 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.815 0.56 4.005 2.475 ;
        RECT 3.815 0.56 4.2 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.37 2.73 2.35 2.92 ;
      RECT 2.115 0.595 2.305 1.31 ;
      RECT 3.39 1.03 3.58 1.31 ;
      RECT 1.265 1.12 3.58 1.31 ;
      RECT 1.265 1.12 1.455 2.475 ;
  END
END AO12V2_7TV50

MACRO AO21BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21BV1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.56 1.32 1.265 ;
        RECT 0.75 1.075 1.32 1.265 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.075 1.97 1.395 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.295 1.04 3.745 1.36 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 2.31 0.505 3.48 ;
        RECT 1.925 2.32 2.205 3.48 ;
        RECT 3.625 2.27 3.905 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.925 -0.12 2.205 0.875 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.82 0.6 3.01 2.475 ;
        RECT 2.82 0.6 3.905 0.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.27 0.595 0.46 1.995 ;
      RECT 0.27 1.805 2.58 1.995 ;
      RECT 1.12 1.805 1.31 2.475 ;
  END
END AO21BV1_7TV50

MACRO AO21BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21BV2_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.72 0.84 2.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.47 1.85 1.86 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.17 1.56 3.76 1.805 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.255 0.39 3.48 ;
        RECT 1.855 2.255 2.135 3.48 ;
        RECT 3.555 2.65 3.835 3.48 ;
        RECT 5.3 2.29 5.535 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.855 -0.12 2.135 0.76 ;
        RECT 5.3 -0.12 5.535 0.71 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 0.56 3.72 0.88 ;
        RECT 3.48 0.64 5.1 0.83 ;
        RECT 4.91 0.64 5.1 2.43 ;
        RECT 2.705 2.24 5.1 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.155 0.64 1.24 0.83 ;
      RECT 1.05 1.08 4.71 1.27 ;
      RECT 4.52 1.08 4.71 1.63 ;
      RECT 1.05 0.64 1.24 2.475 ;
  END
END AO21BV2_7TV50

MACRO AO221V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.775 0.6 3.965 1.31 ;
        RECT 3.775 0.6 4.24 0.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.89 1.36 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.03 2.945 1.34 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.6 2.19 1.31 ;
        RECT 2 0.6 2.32 0.84 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.075 1.46 1.42 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.195 2.63 3.475 3.48 ;
        RECT 4.955 2.295 5.235 3.48 ;
        RECT 3.195 3.215 5.235 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.505 -0.12 1.785 0.835 ;
        RECT 4.905 -0.12 5.185 0.84 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.85 0.56 6.04 2.475 ;
        RECT 5.85 0.56 6.12 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.86 2.24 4.385 2.43 ;
      RECT 3.25 0.59 3.44 1.855 ;
      RECT 0.65 1.665 5.61 1.855 ;
      RECT 0.65 0.595 0.84 2.43 ;
      RECT 0.205 2.24 0.84 2.43 ;
  END
END AO221V1_7TV50

MACRO AO221V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221V2_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.815 0.6 4.005 1.31 ;
        RECT 3.815 0.6 4.24 0.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.89 1.36 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 1.04 2.97 1.36 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.6 2.19 1.31 ;
        RECT 2 0.6 2.32 0.84 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.04 1.5 1.385 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.295 2.645 3.575 3.48 ;
        RECT 4.995 2.255 5.275 3.48 ;
        RECT 6.695 2.275 6.975 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.545 -0.12 1.78 0.795 ;
        RECT 4.945 -0.12 5.225 0.795 ;
        RECT 6.745 -0.12 7.025 0.75 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.89 0.56 6.08 2.475 ;
        RECT 5.88 0.56 6.12 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.75 2.985 2.94 ;
      RECT 1.855 2.24 4.425 2.43 ;
      RECT 0.69 0.595 0.88 1.995 ;
      RECT 3.29 0.59 3.48 1.995 ;
      RECT 0.2 1.805 5.65 1.995 ;
      RECT 0.2 1.805 0.39 2.475 ;
  END
END AO221V2_7TV50

MACRO AO222V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222V1_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.72 0.6 4.91 1.31 ;
        RECT 4.72 0.6 5.2 0.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.29 1.04 5.74 1.36 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.43 0.6 2.62 1.31 ;
        RECT 2.43 0.6 2.8 0.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.995 1.04 3.445 1.36 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.075 1.61 1.33 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.895 2.04 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.2 2.63 4.48 3.48 ;
        RECT 5.9 2.53 6.18 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.875 ;
        RECT 3.56 -0.12 3.84 0.875 ;
        RECT 5.85 -0.12 6.13 0.87 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.795 0.56 6.985 2.475 ;
        RECT 6.795 0.56 7.08 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.255 2.355 0.445 3.02 ;
      RECT 1.955 2.355 2.145 3.02 ;
      RECT 3.655 2.355 3.845 3.02 ;
      RECT 0.255 2.83 3.845 3.02 ;
      RECT 2.805 1.95 5.285 2.14 ;
      RECT 2.805 1.95 2.995 2.475 ;
      RECT 5.095 1.95 5.285 2.705 ;
      RECT 1.905 0.595 2.095 1.75 ;
      RECT 4.195 0.595 4.385 1.75 ;
      RECT 1.105 1.56 6.51 1.75 ;
      RECT 6.32 1.56 6.51 1.94 ;
      RECT 1.105 1.56 1.295 2.475 ;
  END
END AO222V1_7TV50

MACRO AO222V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.665 0.6 4.855 1.31 ;
        RECT 4.665 0.6 5.2 0.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.04 5.85 1.36 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 0.97 3.85 1.36 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 0.6 3.15 1.31 ;
        RECT 2.96 0.6 3.28 0.84 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.52 0.84 2.04 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.865 1.01 2.32 1.33 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.145 2.685 4.425 3.48 ;
        RECT 5.845 2.245 6.125 3.48 ;
        RECT 7.545 2.275 7.825 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.39 -0.12 2.67 0.765 ;
        RECT 5.795 -0.12 6.075 0.76 ;
        RECT 7.595 -0.12 7.875 0.75 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.74 0.56 6.93 2.475 ;
        RECT 6.74 0.56 7.08 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.155 2.73 3.835 2.92 ;
      RECT 2.705 2.24 5.275 2.43 ;
      RECT 0.69 0.64 1.24 0.83 ;
      RECT 4.14 0.595 4.33 1.895 ;
      RECT 1.05 1.705 6.5 1.895 ;
      RECT 1.05 0.64 1.24 2.475 ;
  END
END AO222V2_7TV50

MACRO AO22V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22V1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 1.56 1.84 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.435 1.075 0.88 1.4 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.04 2.515 1.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3 1.52 3.72 1.865 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.09 2.4 1.37 3.48 ;
        RECT 4.23 2.275 4.51 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.19 -0.12 0.47 0.875 ;
        RECT 0.19 -0.12 3.87 0.145 ;
        RECT 3.59 -0.12 3.87 0.875 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.49 0.6 5.315 0.84 ;
        RECT 5.125 0.6 5.315 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.285 2.01 2.175 2.2 ;
      RECT 0.285 2.01 0.475 2.475 ;
      RECT 1.985 2.01 2.175 2.82 ;
      RECT 3.685 2.355 3.875 2.82 ;
      RECT 1.985 2.63 3.875 2.82 ;
      RECT 1.89 0.64 3.025 0.83 ;
      RECT 2.835 1.075 4.245 1.265 ;
      RECT 2.835 0.64 3.025 2.43 ;
      RECT 2.79 2.24 3.07 2.43 ;
  END
END AO22V1_7TV50

MACRO AO22V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22V2_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.245 1.56 1.845 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.555 1.075 1 1.4 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.04 2.62 1.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.3 1.52 3.72 1.865 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.09 2.685 1.37 3.48 ;
        RECT 4.23 2.275 4.51 3.48 ;
        RECT 5.93 2.275 6.21 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.31 -0.12 0.59 0.78 ;
        RECT 0.31 -0.12 3.99 0.145 ;
        RECT 3.71 -0.12 3.99 0.78 ;
        RECT 5.555 -0.12 5.79 0.735 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.61 0.6 5.315 0.84 ;
        RECT 5.125 0.6 5.315 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.24 2.24 2.175 2.43 ;
      RECT 1.985 2.24 2.175 2.92 ;
      RECT 1.985 2.73 3.92 2.92 ;
      RECT 2.01 0.64 3.025 0.83 ;
      RECT 2.835 1.075 4.365 1.265 ;
      RECT 2.835 0.64 3.025 2.475 ;
  END
END AO22V2_7TV50

MACRO AO31V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 0.56 1.8 0.88 ;
        RECT 1.61 0.56 1.8 1.31 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.21 1.075 2.8 1.32 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 0.6 3.28 0.84 ;
        RECT 3.09 0.6 3.28 1.31 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.29 1.075 0.88 1.32 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.905 2.4 2.185 3.48 ;
        RECT 3.605 2.29 3.885 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.875 ;
        RECT 3.555 -0.12 3.835 0.875 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 0.56 4.69 0.88 ;
        RECT 4.5 0.56 4.69 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.1 2.01 2.99 2.2 ;
      RECT 1.1 2.01 1.29 2.475 ;
      RECT 2.8 2.01 2.99 2.475 ;
      RECT 1.1 0.595 1.29 1.765 ;
      RECT 0.25 1.575 4.26 1.765 ;
      RECT 0.25 1.575 0.44 2.475 ;
  END
END AO31V1_7TV50

MACRO AO31V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 0.56 1.8 0.88 ;
        RECT 1.61 0.56 1.8 1.31 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.38 1.075 2.8 1.42 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 0.6 3.28 0.84 ;
        RECT 3.09 0.6 3.28 1.31 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.53 1.06 0.88 1.475 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.905 2.685 2.185 3.48 ;
        RECT 3.605 2.29 3.885 3.48 ;
        RECT 5.305 2.28 5.585 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.86 ;
        RECT 3.555 -0.12 3.835 0.79 ;
        RECT 5.355 -0.12 5.635 0.745 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 0.495 4.69 0.88 ;
        RECT 4.5 0.495 4.69 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.055 2.24 3.035 2.43 ;
      RECT 1.1 0.595 1.29 1.945 ;
      RECT 0.25 1.755 4.26 1.945 ;
      RECT 0.25 1.755 0.44 2.475 ;
  END
END AO31V2_7TV50

MACRO AO32V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32V1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.315 1.485 2.81 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.98 1.04 3.495 1.365 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.92 1.485 4.385 1.84 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5 1.02 1.97 1.37 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.44 1.52 0.89 1.9 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.705 2.4 2.985 3.48 ;
        RECT 4.405 2.4 4.685 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.82 ;
        RECT 4.355 -0.12 4.635 0.82 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.3 0.57 5.49 2.475 ;
        RECT 5.3 1.52 5.64 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.9 2.01 3.72 2.2 ;
      RECT 3.53 2.01 3.72 2.585 ;
      RECT 3.53 2.395 3.835 2.585 ;
      RECT 0.2 2.355 0.39 2.985 ;
      RECT 1.9 2.01 2.09 2.985 ;
      RECT 0.2 2.795 2.09 2.985 ;
      RECT 1.09 0.63 4.155 0.82 ;
      RECT 3.965 0.63 4.155 1.255 ;
      RECT 3.965 1.065 5.01 1.255 ;
      RECT 1.09 0.63 1.29 2.59 ;
      RECT 1.005 2.4 1.29 2.59 ;
  END
END AO32V1_7TV50

MACRO AO32V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32V2_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.36 1.49 2.76 1.94 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.22 1.065 3.77 1.375 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.075 1.51 4.68 1.85 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.51 1.03 1.975 1.38 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.455 1.49 0.85 1.94 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.79 2.73 3.07 3.48 ;
        RECT 4.49 2.34 4.77 3.48 ;
        RECT 6.19 2.4 6.47 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 -0.12 0.485 0.66 ;
        RECT 4.405 -0.12 4.685 0.66 ;
        RECT 6.205 -0.12 6.485 0.58 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.35 0.595 5.54 2.43 ;
        RECT 5.34 2.24 5.62 2.43 ;
        RECT 5.35 1.04 5.64 1.36 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.17 2.295 3.92 2.485 ;
      RECT 2.17 2.295 2.36 2.82 ;
      RECT 0.24 2.63 2.36 2.82 ;
      RECT 1.12 0.64 4.205 0.83 ;
      RECT 4.015 0.64 4.205 1.22 ;
      RECT 4.015 1.03 5.015 1.22 ;
      RECT 4.825 1.03 5.015 1.31 ;
      RECT 1.12 0.64 1.31 2.43 ;
      RECT 1.09 2.24 1.37 2.43 ;
  END
END AO32V2_7TV50

MACRO AO33V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.08 3.405 1.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.805 1.08 4.255 1.4 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.92 1.52 5.25 1.98 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.52 2.555 1.85 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.475 1.08 1.84 1.475 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.42 1.03 0.84 1.405 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.6 2.4 3.88 3.48 ;
        RECT 5.3 2.4 5.58 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.2 -0.12 0.48 0.815 ;
        RECT 5.25 -0.12 5.53 0.815 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.195 0.56 6.385 2.475 ;
        RECT 6.195 1.52 6.6 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.795 1.965 4.685 2.155 ;
      RECT 4.495 1.965 4.685 2.475 ;
      RECT 1.095 2.355 1.285 2.82 ;
      RECT 2.795 1.965 2.99 2.82 ;
      RECT 1.095 2.63 2.99 2.82 ;
      RECT 1.085 0.625 4.77 0.815 ;
      RECT 4.58 0.625 4.77 1.25 ;
      RECT 4.58 1.06 5.905 1.25 ;
      RECT 1.085 0.625 1.275 2.055 ;
      RECT 0.245 1.865 1.675 2.055 ;
      RECT 1.485 1.865 1.675 2.43 ;
      RECT 1.485 2.24 2.18 2.43 ;
      RECT 0.245 1.865 0.435 2.475 ;
  END
END AO33V1_7TV50

MACRO AO33V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33V2_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.525 1.95 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.895 1 4.345 1.32 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.88 1.445 5.26 1.825 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.56 2.595 1.95 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 0.99 1.95 1.36 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 1.52 0.895 1.845 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.69 2.73 3.97 3.48 ;
        RECT 5.515 2.34 5.795 3.48 ;
        RECT 7.215 2.4 7.495 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.19 -0.12 0.47 0.66 ;
        RECT 5.415 -0.12 5.695 0.66 ;
        RECT 7.215 -0.12 7.495 0.58 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.315 0.56 6.6 0.75 ;
        RECT 6.36 1.52 6.6 1.84 ;
        RECT 6.41 0.56 6.6 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.07 2.34 4.82 2.53 ;
      RECT 3.07 2.34 3.26 2.82 ;
      RECT 1.09 2.63 3.26 2.82 ;
      RECT 1.17 0.56 5.215 0.75 ;
      RECT 5.025 0.56 5.215 1.05 ;
      RECT 5.025 0.86 6.13 1.05 ;
      RECT 5.94 0.86 6.13 1.31 ;
      RECT 1.17 0.56 1.36 2.43 ;
      RECT 0.24 2.24 2.22 2.43 ;
  END
END AO33V2_7TV50

MACRO AOI211V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.52 1.81 1.985 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 1.01 0.915 1.36 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.325 1.5 2.8 1.855 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.94 1.265 4.22 1.84 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 2.79 1.335 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.58 ;
        RECT 2.755 -0.12 3.035 0.58 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.9 0.595 2.09 0.97 ;
        RECT 3.48 1.995 3.74 2.32 ;
        RECT 3.55 0.78 3.74 2.475 ;
        RECT 3.7 0.595 3.89 0.97 ;
        RECT 1.9 0.78 3.89 0.97 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.205 2.24 2.185 2.43 ;
  END
END AOI211V1_7TV50

MACRO AOI211V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.51 1.08 1.86 1.32 ;
        RECT 1.51 1.08 2.76 1.27 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 0.88 1.8 ;
        RECT 0.56 1.61 3.365 1.8 ;
        RECT 3.175 1.61 3.365 2.04 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4 1.08 4.72 1.32 ;
        RECT 4.15 1.08 6.385 1.27 ;
        RECT 6.195 1.08 6.385 1.6 ;
        RECT 6.195 1.41 6.64 1.6 ;
        RECT 6.45 1.41 6.64 2.04 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.52 5.64 1.995 ;
        RECT 4.83 1.805 5.96 1.995 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 2.79 1.335 3.48 ;
        RECT 2.755 2.79 3.035 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 -0.12 0.535 0.58 ;
        RECT 3.715 -0.12 3.995 0.39 ;
        RECT 5.635 -0.12 5.915 0.39 ;
        RECT 7.495 -0.12 7.775 0.58 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.955 0.64 7.03 0.83 ;
        RECT 6.84 0.64 7.03 2.43 ;
        RECT 5.205 2.24 7.03 2.43 ;
        RECT 6.84 1.52 7.08 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.19 2.24 3.655 2.43 ;
      RECT 3.465 2.24 3.655 2.98 ;
      RECT 3.465 2.79 7.225 2.98 ;
  END
END AOI211V2_7TV50

MACRO AOI21BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BV1_7TV50 0 0 ;
  SIZE 4.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.12 1.485 0.53 1.84 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.885 1.04 3.26 1.425 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.8 1.52 4.2 1.88 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 2.365 1.315 3.48 ;
        RECT 3.37 2.79 3.65 3.48 ;
        RECT 0 3.24 4.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.56 -0.12 1.84 0.39 ;
        RECT 4.22 -0.12 4.5 0.58 ;
        RECT 0 -0.12 4.8 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.715 0.65 1.905 2.475 ;
        RECT 2.48 0.6 2.8 0.84 ;
        RECT 1.715 0.65 2.8 0.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.18 0.64 1.51 0.83 ;
      RECT 1.32 0.64 1.51 1.82 ;
      RECT 0.73 1.63 1.51 1.82 ;
      RECT 0.73 1.63 0.92 2.385 ;
      RECT 0.275 2.195 0.92 2.385 ;
      RECT 0.275 2.195 0.465 2.475 ;
      RECT 2.52 2.24 4.5 2.43 ;
  END
END AOI21BV1_7TV50

MACRO AOI21BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21BV2_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.495 1.765 0.84 2.32 ;
        RECT 0.415 2 0.84 2.32 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.36 1.08 5.68 1.41 ;
        RECT 4.255 1.22 5.68 1.41 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.735 1.61 4.055 2.005 ;
        RECT 6.365 1.56 6.56 2.05 ;
        RECT 6.32 1.56 6.64 1.8 ;
        RECT 3.735 1.61 6.64 1.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.635 0.435 3.48 ;
        RECT 4.145 2.795 4.425 3.48 ;
        RECT 5.845 2.795 6.125 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.565 ;
        RECT 2.855 -0.12 3.135 0.565 ;
        RECT 6.575 -0.12 6.855 0.565 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.58 2.19 0.99 ;
        RECT 2.49 0.8 2.68 2.485 ;
        RECT 2.49 1.52 2.76 1.84 ;
        RECT 4.715 0.71 4.995 0.99 ;
        RECT 2 0.8 4.995 0.99 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.2 -0.24 5.345 1.53 ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.2 3.94 ;
        RECT 5.345 1.46 7.78 3.94 ;
        RECT -0.58 1.53 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 0.5 0.39 1.325 ;
      RECT 0.2 1.135 1.86 1.325 ;
      RECT 1.05 1.135 1.24 2.48 ;
      RECT 3.755 0.32 5.955 0.51 ;
      RECT 3.755 0.32 4.035 0.565 ;
      RECT 5.675 0.32 5.955 0.565 ;
      RECT 3.155 2.405 6.975 2.595 ;
      RECT 3.155 2.405 3.345 2.985 ;
      RECT 1.595 2.795 3.345 2.985 ;
  END
END AOI21BV2_7TV50

MACRO AOI21V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.33 1.46 2.8 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.45 1.945 1.8 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.74 0.85 2.32 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.855 2.79 2.135 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.58 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2 0.59 0.39 2.475 ;
        RECT 2.52 0.56 3.035 0.97 ;
        RECT 0.2 0.78 3.035 0.97 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.05 2.24 2.985 2.43 ;
      RECT 1.05 2.24 1.24 2.78 ;
  END
END AOI21V1_7TV50

MACRO AOI21V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.74 1.08 4.285 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.56 2.8 1.8 ;
        RECT 2.48 1.61 5.2 1.8 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.42 1.005 0.88 1.32 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.855 2.79 3.135 3.48 ;
        RECT 4.655 2.79 4.935 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 -0.12 0.485 0.625 ;
        RECT 2.005 -0.12 2.285 0.58 ;
        RECT 5.455 -0.12 5.735 0.625 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.52 1.34 1.84 ;
        RECT 1.15 0.515 1.34 2.475 ;
        RECT 1.15 0.825 3.17 1.025 ;
        RECT 2.93 0.64 4.035 0.83 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.05 2.4 5.785 2.59 ;
      RECT 2.05 2.4 2.24 2.865 ;
      RECT 0.255 2.675 2.24 2.865 ;
  END
END AOI21V2_7TV50

MACRO AOI221V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221V1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.465 1.945 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 1.065 1.365 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.41 1.47 2.8 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.375 1.42 3.72 1.84 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.41 4.775 1.84 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.25 2.745 1.53 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.4 -0.12 0.68 0.625 ;
        RECT 3.86 -0.12 4.14 0.58 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.145 0.595 2.335 0.97 ;
        RECT 4.865 0.595 5.055 0.97 ;
        RECT 2.145 0.78 5.485 0.97 ;
        RECT 5.295 0.78 5.485 2.475 ;
        RECT 5.295 1.52 5.64 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.4 2.24 4.08 2.43 ;
      RECT 2.95 2.75 4.67 2.94 ;
  END
END AOI221V1_7TV50

MACRO AOI221V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221V2_7TV50 0 0 ;
  SIZE 10.08 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.23 1.08 8.785 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.24 1.52 9.48 1.84 ;
        RECT 6.815 1.65 9.48 1.84 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.91 1.04 4.325 1.31 ;
        RECT 3.96 1.04 4.325 1.41 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.88 1.56 5.235 1.8 ;
        RECT 2.57 1.61 5.235 1.8 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.515 1.495 0.845 1.95 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 6.17 2.745 6.45 3.48 ;
        RECT 7.87 2.745 8.15 3.48 ;
        RECT 9.57 2.355 9.85 3.48 ;
        RECT 0 3.24 10.08 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.12 0.445 0.625 ;
        RECT 1.965 -0.12 2.245 0.625 ;
        RECT 5.785 -0.12 6.455 0.58 ;
        RECT 5.785 -0.12 9.9 0.135 ;
        RECT 9.62 -0.12 9.9 0.625 ;
        RECT 0 -0.12 10.08 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.065 0.595 1.255 2.475 ;
        RECT 1.065 0.595 1.3 1.015 ;
        RECT 1.065 0.825 3.05 1.015 ;
        RECT 2.86 0.6 3.28 0.84 ;
        RECT 2.86 0.64 4.705 0.84 ;
        RECT 4.515 0.78 7.31 0.97 ;
        RECT 7.12 0.64 8.2 0.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 10.2 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 10.66 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.155 2.79 5.695 2.98 ;
      RECT 2.765 2.24 9 2.43 ;
  END
END AOI221V2_7TV50

MACRO AOI222V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.77 1.56 5.2 1.93 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.79 1.56 6.185 1.935 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.845 1.56 4.24 1.94 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.355 1.94 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5 1.52 1.8 2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.42 1.03 0.86 1.36 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.3 2.355 0.58 3.48 ;
        RECT 2 2.76 2.28 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.25 -0.12 0.53 0.62 ;
        RECT 2.64 -0.12 2.92 0.62 ;
        RECT 6.12 -0.12 6.4 0.7 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 0.59 2.23 1.27 ;
        RECT 3.44 1.08 3.76 1.32 ;
        RECT 4.445 0.59 4.635 1.27 ;
        RECT 2.04 1.08 5.59 1.27 ;
        RECT 5.4 1.08 5.59 2.43 ;
        RECT 5.27 2.24 5.59 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.15 2.24 3.83 2.43 ;
      RECT 2.7 2.79 6.415 2.98 ;
  END
END AOI222V1_7TV50

MACRO AOI222V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222V2_7TV50 0 0 ;
  SIZE 11.52 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.28 1.08 1.84 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 0.885 1.8 ;
        RECT 0.56 1.56 3.235 1.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.785 1.08 5.305 1.36 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4 1.56 4.72 1.8 ;
        RECT 4.105 1.61 6.685 1.8 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.645 1.56 10.245 1.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.145 1.115 10.96 1.305 ;
        RECT 10.64 1.08 10.96 1.32 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 8.52 2.79 8.8 3.48 ;
        RECT 10.22 2.79 10.5 3.48 ;
        RECT 0 3.24 11.52 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.275 -0.12 0.465 0.625 ;
        RECT 3.63 -0.12 3.91 0.58 ;
        RECT 7.25 -0.12 7.53 0.58 ;
        RECT 11.02 -0.12 11.3 0.625 ;
        RECT 0 -0.12 11.52 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.93 0.6 3.015 0.84 ;
        RECT 3.655 0.78 3.845 2.445 ;
        RECT 1.08 2.255 3.845 2.445 ;
        RECT 2.825 0.78 4.54 0.97 ;
        RECT 4.35 0.64 6.405 0.83 ;
        RECT 6.215 0.825 7.92 1.015 ;
        RECT 7.73 0.6 9.6 0.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 11.64 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 12.1 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.23 2.79 7.36 2.98 ;
      RECT 4.53 2.24 11.35 2.43 ;
  END
END AOI222V2_7TV50

MACRO AOI22BBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22BBV1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 1.075 0.91 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.54 1.465 1.9 1.865 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.515 3.525 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.285 1.52 4.735 1.84 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.025 2.355 2.305 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.12 0.445 0.875 ;
        RECT 2.025 -0.12 2.32 0.625 ;
        RECT 4.645 -0.12 4.925 0.625 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.925 0.6 4 0.79 ;
        RECT 3.44 0.6 4 0.84 ;
        RECT 3.81 0.6 4 2.475 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.11 1.075 2.68 1.265 ;
      RECT 1.11 0.595 1.3 2.43 ;
      RECT 0.31 2.24 1.3 2.43 ;
      RECT 2.915 2.79 4.895 2.98 ;
  END
END AOI22BBV1_7TV50

MACRO AOI22BBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22BBV2_7TV50 0 0 ;
  SIZE 8.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 1.075 0.91 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.54 1.465 1.9 1.865 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.805 1.555 6.385 1.805 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.67 1.555 8.27 1.805 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.025 2.35 2.305 3.48 ;
        RECT 3.775 2.785 4.055 3.48 ;
        RECT 0 3.24 8.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.12 0.445 0.705 ;
        RECT 2.025 -0.12 2.32 0.625 ;
        RECT 3.825 -0.12 4.105 0.625 ;
        RECT 7.285 -0.12 7.565 0.57 ;
        RECT 0 -0.12 8.64 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.97 0.555 3.16 1.27 ;
        RECT 3.92 1.08 4.24 1.32 ;
        RECT 4.65 1.08 4.84 2.545 ;
        RECT 5.375 0.71 5.655 1.27 ;
        RECT 2.97 1.08 5.655 1.27 ;
        RECT 4.65 2.355 8.465 2.545 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 5.07 -0.24 5.96 1.53 ;
        RECT -0.12 -0.24 8.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.07 3.94 ;
        RECT 5.96 1.46 9.22 3.94 ;
        RECT -0.58 1.53 9.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.11 1.075 2.68 1.265 ;
      RECT 1.11 0.595 1.3 2.43 ;
      RECT 0.315 2.24 1.3 2.43 ;
      RECT 2.875 2.395 4.445 2.585 ;
      RECT 4.255 2.395 4.445 2.985 ;
      RECT 4.255 2.795 7.565 2.985 ;
      RECT 4.46 0.32 6.615 0.51 ;
      RECT 4.46 0.32 4.65 0.615 ;
      RECT 6.425 0.32 6.615 0.97 ;
      RECT 8.23 0.585 8.42 0.97 ;
      RECT 6.425 0.77 8.42 0.97 ;
  END
END AOI22BBV2_7TV50

MACRO AOI22V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.545 1.52 1.86 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5 1.55 1.01 1.815 ;
        RECT 0.73 1.55 1.01 1.995 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.36 1.03 2.76 1.39 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.425 1.505 3.76 1.995 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.79 1.485 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.355 -0.12 0.635 0.625 ;
        RECT 3.755 -0.12 4.035 0.625 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.055 0.64 3.19 0.83 ;
        RECT 3 0.64 3.19 2.475 ;
        RECT 3 1.04 3.24 1.36 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.355 2.24 2.525 2.43 ;
      RECT 2.335 2.24 2.525 2.865 ;
      RECT 2.335 2.675 4.085 2.865 ;
  END
END AOI22V1_7TV50

MACRO AOI22V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.84 1.08 6.33 1.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4 1.56 4.72 1.8 ;
        RECT 4.4 1.61 7.26 1.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.895 1.08 2.325 1.32 ;
        RECT 1.895 1.08 2.925 1.27 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.515 1.56 1.84 1.8 ;
        RECT 1.095 1.61 3.76 1.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.87 2.75 5.15 3.48 ;
        RECT 6.575 2.75 6.855 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.57 -0.12 0.85 0.595 ;
        RECT 3.97 -0.12 4.25 0.58 ;
        RECT 7.375 -0.12 7.655 0.625 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.27 0.64 3.39 0.83 ;
        RECT 3.96 2 4.2 2.43 ;
        RECT 4.01 0.78 4.2 2.43 ;
        RECT 1.37 2.24 4.2 2.43 ;
        RECT 3.2 0.78 5.545 0.97 ;
        RECT 5.355 0.64 5.95 0.83 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 4.45 2.355 7.705 2.545 ;
      RECT 4.45 2.355 4.64 2.82 ;
      RECT 0.52 2.63 4.64 2.82 ;
  END
END AOI22V2_7TV50

MACRO AOI22XBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22XBV1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.41 1.465 1.84 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.355 1.54 0.91 1.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.04 2.53 1.36 ;
    END
  END B1
  PIN B2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.39 1.465 4.715 1.91 ;
    END
  END B2N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.02 2.79 1.3 3.48 ;
        RECT 4.16 2.205 4.44 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.17 -0.12 0.45 0.65 ;
        RECT 3.57 -0.12 3.85 0.65 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.87 0.6 2.955 0.79 ;
        RECT 2.48 0.6 2.955 0.84 ;
        RECT 2.765 0.6 2.955 2.475 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.17 2.4 2.105 2.59 ;
      RECT 1.915 2.4 2.105 2.865 ;
      RECT 1.915 2.675 3.85 2.865 ;
      RECT 4.575 0.595 4.765 1.265 ;
      RECT 3.195 1.075 5.245 1.265 ;
      RECT 5.055 1.075 5.245 2.485 ;
  END
END AOI22XBV1_7TV50

MACRO AOI22XBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22XBV2_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.46 1.04 8.04 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.665 1.56 6.18 1.81 ;
        RECT 5.665 1.62 8.285 1.81 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.755 1.08 3.295 1.35 ;
    END
  END B1
  PIN B2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.08 0.955 1.335 ;
    END
  END B2N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.3 2.41 0.58 3.48 ;
        RECT 6.04 2.79 6.32 3.48 ;
        RECT 7.79 2.79 8.07 3.48 ;
        RECT 6.04 3.235 8.07 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 -0.12 0.485 0.745 ;
        RECT 1.79 -0.12 2.07 0.625 ;
        RECT 5.19 -0.12 5.47 0.625 ;
        RECT 1.79 -0.12 8.87 0.135 ;
        RECT 8.59 -0.12 8.87 0.625 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.535 0.595 3.725 1.275 ;
        RECT 4.4 1.08 4.72 1.32 ;
        RECT 5.26 1.08 5.45 2.43 ;
        RECT 2.59 2.24 5.45 2.43 ;
        RECT 6.935 0.595 7.125 1.275 ;
        RECT 3.535 1.08 7.125 1.275 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.195 1.805 4.995 1.995 ;
      RECT 1.195 0.595 1.385 2.475 ;
      RECT 5.65 2.4 8.92 2.59 ;
      RECT 5.65 2.4 5.84 2.86 ;
      RECT 1.74 2.67 5.84 2.86 ;
  END
END AOI22XBV2_7TV50

MACRO AOI2XB11V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB11V1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.995 1.56 2.595 1.8 ;
    END
  END A1
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.49 1.425 0.84 1.84 ;
    END
  END A2N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.285 1.56 3.945 1.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.78 1.56 5.38 1.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.205 0.435 3.48 ;
        RECT 2.585 2.79 2.865 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.685 -0.12 1.965 0.83 ;
        RECT 4.345 -0.12 4.625 0.74 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.43 0.58 3.62 1.27 ;
        RECT 3.915 1.08 4.51 1.32 ;
        RECT 4.32 1.08 4.51 2.43 ;
        RECT 4.32 2.24 5.315 2.43 ;
        RECT 5.35 0.595 5.54 1.27 ;
        RECT 3.43 1.08 5.54 1.27 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.75 0.64 1.24 0.83 ;
      RECT 1.04 1.075 3.14 1.265 ;
      RECT 1.04 0.64 1.24 2.475 ;
      RECT 1.735 2.24 3.715 2.43 ;
  END
END AOI2XB11V1_7TV50

MACRO AOI2XB11V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB11V2_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.56 3.76 1.8 ;
        RECT 2.09 1.61 4.75 1.8 ;
    END
  END A1
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.415 1.865 0.84 2.115 ;
        RECT 0.6 1.865 0.84 2.32 ;
    END
  END A2N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.74 1.08 8.08 1.345 ;
        RECT 5.48 1.08 8.44 1.27 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.515 1.56 7.12 1.825 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 2.665 0.455 3.48 ;
        RECT 2.465 2.79 2.745 3.48 ;
        RECT 4.27 2.79 4.55 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.445 -0.12 1.725 0.745 ;
        RECT 4.905 -0.12 5.185 0.44 ;
        RECT 6.825 -0.12 7.105 0.44 ;
        RECT 8.685 -0.12 8.965 0.625 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.92 0.64 5.16 1.36 ;
        RECT 4.97 0.64 5.16 1.8 ;
        RECT 4.97 1.61 6.07 1.8 ;
        RECT 5.88 1.61 6.07 2.43 ;
        RECT 5.88 2.24 7.205 2.43 ;
        RECT 3.145 0.64 8.065 0.83 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.59 0.595 0.78 1.34 ;
      RECT 0.59 1.15 2.92 1.34 ;
      RECT 1.07 1.15 1.26 2.565 ;
      RECT 1.615 2.24 5.355 2.43 ;
      RECT 5.165 2.24 5.355 2.865 ;
      RECT 5.165 2.675 8.825 2.865 ;
  END
END AOI2XB11V2_7TV50

MACRO AOI2XB1V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1V1_7TV50 0 0 ;
  SIZE 4.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.94 1.04 4.68 1.29 ;
        RECT 4.44 1.04 4.68 1.36 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.965 3.24 1.565 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.495 1.56 0.93 1.895 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 2.195 0.495 3.48 ;
        RECT 2.615 2.79 2.895 3.48 ;
        RECT 0 3.24 4.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.875 ;
        RECT 1.715 -0.12 1.995 0.625 ;
        RECT 1.715 -0.12 4.595 0.135 ;
        RECT 4.3 -0.12 4.595 0.625 ;
        RECT 0 -0.12 4.8 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.46 0.595 3.65 1.75 ;
        RECT 3.46 1.56 4.55 1.75 ;
        RECT 3.92 1.56 4.55 1.8 ;
        RECT 4.36 1.56 4.55 2.475 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.17 1.075 2.37 1.265 ;
      RECT 1.17 0.595 1.36 2.475 ;
      RECT 1.765 2.24 3.745 2.43 ;
  END
END AOI2XB1V1_7TV50

MACRO AOI2XB1V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2XB1V2_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.36 1.04 6.81 1.36 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.68 1.08 3.28 1.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.495 1.04 0.955 1.36 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.26 2.195 0.54 3.48 ;
        RECT 2.565 2.79 2.845 3.48 ;
        RECT 4.265 2.79 4.545 3.48 ;
        RECT 2.565 3.235 4.545 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.21 -0.12 0.49 0.745 ;
        RECT 1.765 -0.12 2.045 0.625 ;
        RECT 5.165 -0.12 5.445 0.625 ;
        RECT 6.965 -0.12 7.245 0.625 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.51 0.595 3.7 1.27 ;
        RECT 4.88 1.08 5.2 1.32 ;
        RECT 3.51 1.08 6.16 1.27 ;
        RECT 5.97 0.64 6.16 2.475 ;
        RECT 5.97 2.195 6.2 2.475 ;
        RECT 5.97 0.64 6.345 0.83 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.11 0.64 1.39 0.83 ;
      RECT 1.2 1.575 4.92 1.765 ;
      RECT 1.2 0.64 1.39 2.43 ;
      RECT 1.11 2.24 1.39 2.43 ;
      RECT 1.7 2.24 5.35 2.43 ;
      RECT 5.16 2.24 5.35 2.865 ;
      RECT 5.16 2.675 7.095 2.865 ;
  END
END AOI2XB1V2_7TV50

MACRO AOI31V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.56 2.465 1.87 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.385 1.01 1.8 1.36 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.415 1.5 0.84 1.84 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.18 1.07 3.76 1.32 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.27 0.435 3.48 ;
        RECT 1.855 2.665 2.135 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.73 ;
        RECT 3.555 -0.12 3.835 0.7 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.7 0.595 2.89 1.8 ;
        RECT 2.7 1.56 3.79 1.8 ;
        RECT 3.6 1.56 3.79 2.475 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.275 2.985 2.465 ;
  END
END AOI31V1_7TV50

MACRO AOI31V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31V2_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.6 2.42 0.84 ;
        RECT 2.23 0.6 2.42 1.125 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.525 1.04 1.8 1.515 ;
        RECT 1.525 1.325 4.22 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.84 1.905 ;
        RECT 0.6 1.715 5.12 1.905 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.64 1.515 7.15 1.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.695 1.345 3.48 ;
        RECT 2.765 2.695 3.045 3.48 ;
        RECT 4.465 2.695 4.745 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.75 ;
        RECT 5.265 -0.12 5.545 0.75 ;
        RECT 7.065 -0.12 7.345 0.75 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.71 0.455 4.63 0.645 ;
        RECT 4.44 0.455 4.63 1.36 ;
        RECT 4.44 1.04 4.68 1.36 ;
        RECT 4.44 1.17 6.4 1.36 ;
        RECT 6.21 0.595 6.4 2.48 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.215 2.245 5.55 2.435 ;
      RECT 5.36 2.245 5.55 2.985 ;
      RECT 5.36 2.795 7.295 2.985 ;
  END
END AOI31V2_7TV50

MACRO AOI32V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 0.915 2.365 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 1.56 1.84 1.81 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.43 1 0.88 1.32 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.385 3.315 1.845 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 1.04 4.41 1.36 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.275 0.435 3.48 ;
        RECT 1.855 2.745 2.135 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.75 ;
        RECT 4.355 -0.12 4.635 0.75 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.655 0.6 3.745 0.84 ;
        RECT 3.555 0.6 3.745 2.43 ;
        RECT 3.555 2.24 3.835 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.355 2.94 2.545 ;
      RECT 2.75 2.355 2.94 2.98 ;
      RECT 2.75 2.79 4.685 2.98 ;
  END
END AOI32V1_7TV50

MACRO AOI32V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32V2_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.6 2.42 0.84 ;
        RECT 2.23 0.6 2.42 1.125 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.525 1.04 1.8 1.515 ;
        RECT 1.525 1.325 4.22 1.515 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.84 1.905 ;
        RECT 0.6 1.715 5.06 1.905 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.49 1.075 8.08 1.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.73 1.56 8.56 1.75 ;
        RECT 8.24 1.56 8.56 1.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.74 1.285 3.48 ;
        RECT 2.705 2.74 2.985 3.48 ;
        RECT 4.405 2.74 4.685 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.75 ;
        RECT 5.265 -0.12 5.545 0.625 ;
        RECT 8.665 -0.12 8.945 0.75 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.755 0.41 2.945 1.07 ;
        RECT 5.3 0.88 5.49 2.14 ;
        RECT 6.15 1.95 6.34 2.48 ;
        RECT 7.01 0.595 7.2 1.07 ;
        RECT 2.755 0.88 7.2 1.07 ;
        RECT 5.3 1.95 8.04 2.14 ;
        RECT 7.8 1.95 8.04 2.48 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.155 2.35 5.49 2.54 ;
      RECT 5.3 2.35 5.49 2.985 ;
      RECT 5.3 2.795 8.935 2.985 ;
  END
END AOI32V2_7TV50

MACRO BUFV16_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV16_7TV50 0 0 ;
  SIZE 20.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.485 3.28 1.8 ;
        RECT 1.795 1.485 4.21 1.675 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.16 2.3 0.44 3.48 ;
        RECT 1.995 2.745 2.275 3.48 ;
        RECT 3.71 2.745 3.99 3.48 ;
        RECT 5.56 2.27 5.84 3.48 ;
        RECT 7.36 2.745 7.64 3.48 ;
        RECT 9.11 2.745 9.39 3.48 ;
        RECT 10.91 2.745 11.19 3.48 ;
        RECT 12.71 2.745 12.99 3.48 ;
        RECT 14.51 2.745 14.79 3.48 ;
        RECT 16.31 2.745 16.59 3.48 ;
        RECT 18.11 2.745 18.39 3.48 ;
        RECT 19.96 2.745 20.24 3.48 ;
        RECT 0 3.24 20.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.16 -0.12 0.44 0.61 ;
        RECT 1.96 -0.12 2.24 0.565 ;
        RECT 3.76 -0.12 4.04 0.565 ;
        RECT 5.56 -0.12 5.84 0.61 ;
        RECT 7.36 -0.12 7.64 0.565 ;
        RECT 9.16 -0.12 9.44 0.565 ;
        RECT 10.96 -0.12 11.24 0.565 ;
        RECT 12.76 -0.12 13.04 0.565 ;
        RECT 14.56 -0.12 14.84 0.565 ;
        RECT 16.36 -0.12 16.64 0.565 ;
        RECT 18.16 -0.12 18.44 0.565 ;
        RECT 19.96 -0.12 20.24 0.61 ;
        RECT 0 -0.12 20.64 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.505 0.595 6.695 0.955 ;
        RECT 8.305 0.595 8.495 0.955 ;
        RECT 10.105 0.595 10.295 0.955 ;
        RECT 11.905 0.595 12.095 0.955 ;
        RECT 12.6 0.765 12.84 1.36 ;
        RECT 12.65 0.765 12.84 2.545 ;
        RECT 13.705 0.595 13.895 0.955 ;
        RECT 15.505 0.595 15.695 0.955 ;
        RECT 17.305 0.595 17.495 0.955 ;
        RECT 19.105 0.595 19.295 0.955 ;
        RECT 6.505 0.765 19.295 0.955 ;
        RECT 6.46 2.355 19.34 2.545 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 20.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 21.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.105 0.595 1.295 0.955 ;
      RECT 2.905 0.595 3.095 0.955 ;
      RECT 1.105 0.765 4.895 0.955 ;
      RECT 4.705 1.485 12.315 1.675 ;
      RECT 4.705 0.595 4.895 2.54 ;
      RECT 1.145 2.35 4.895 2.54 ;
  END
END BUFV16_7TV50

MACRO BUFV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV1_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.91 1.52 1.32 1.875 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 2.75 1.395 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 -0.12 1.345 0.875 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.965 0.64 2.245 0.83 ;
        RECT 2.055 0.64 2.245 2.43 ;
        RECT 1.965 2.24 2.245 2.43 ;
        RECT 2.04 1.52 2.28 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.205 0.595 0.395 2.43 ;
      RECT 1.535 1.76 1.725 2.43 ;
      RECT 0.205 2.24 1.725 2.43 ;
  END
END BUFV1_7TV50

MACRO BUFV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV2_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.925 1.49 1.32 1.855 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.155 2.685 1.435 3.48 ;
        RECT 2.895 2.325 3.175 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.09 -0.12 1.375 0.65 ;
        RECT 2.895 -0.12 3.175 0.695 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 0.575 2.23 3.015 ;
        RECT 2.04 1.52 2.28 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.24 0.595 0.43 2.43 ;
      RECT 1.575 1.76 1.765 2.43 ;
      RECT 0.24 2.24 1.765 2.43 ;
  END
END BUFV2_7TV50

MACRO BUFV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV3_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.75 1.08 0.94 1.36 ;
        RECT 0.75 1.08 1.36 1.32 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.08 2.345 1.36 3.48 ;
        RECT 2.88 2.75 3.16 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.08 -0.12 1.36 0.61 ;
        RECT 2.88 -0.12 3.16 0.565 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.025 0.595 2.215 0.955 ;
        RECT 2.025 0.765 4.015 0.955 ;
        RECT 3.44 2.04 4.015 2.43 ;
        RECT 3.825 0.595 4.015 2.43 ;
        RECT 2.03 2.24 4.015 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.18 0.64 0.465 0.83 ;
      RECT 0.275 1.65 1.885 1.84 ;
      RECT 0.275 0.64 0.465 2.475 ;
  END
END BUFV3_7TV50

MACRO BUFV4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV4_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 1.56 1.375 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.375 2.52 0.655 3.48 ;
        RECT 2.175 2.415 2.455 3.48 ;
        RECT 4.025 2.675 4.305 3.48 ;
        RECT 5.775 2.395 6.055 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.375 -0.12 0.655 0.76 ;
        RECT 2.175 -0.12 2.455 0.76 ;
        RECT 3.975 -0.12 4.255 0.565 ;
        RECT 5.775 -0.12 6.055 0.61 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.12 0.595 3.31 0.955 ;
        RECT 4.875 0.63 5.16 0.955 ;
        RECT 3.12 0.765 5.16 0.955 ;
        RECT 4.92 1.52 5.16 1.84 ;
        RECT 4.97 0.63 5.16 2.43 ;
        RECT 3.175 2.24 5.16 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.275 0.64 1.765 0.83 ;
      RECT 1.575 1.45 3.61 1.64 ;
      RECT 1.575 0.64 1.765 2.55 ;
      RECT 1.325 2.36 1.765 2.55 ;
  END
END BUFV4_7TV50

MACRO BUFV6_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV6_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.83 1.56 1.36 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.36 2.335 0.64 3.48 ;
        RECT 2.205 2.335 2.485 3.48 ;
        RECT 4.01 2.745 4.29 3.48 ;
        RECT 5.755 2.745 6.035 3.48 ;
        RECT 7.605 2.345 7.885 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.36 -0.12 0.64 0.61 ;
        RECT 2.205 -0.12 2.485 0.61 ;
        RECT 4.005 -0.12 4.285 0.565 ;
        RECT 5.805 -0.12 6.085 0.565 ;
        RECT 7.605 -0.12 7.885 0.61 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.15 0.58 3.34 0.955 ;
        RECT 4.95 0.58 5.14 2.43 ;
        RECT 4.92 0.765 5.16 1.36 ;
        RECT 6.75 0.58 6.94 0.955 ;
        RECT 3.15 0.765 6.94 0.955 ;
        RECT 3.135 2.24 6.985 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.305 0.635 1.75 0.835 ;
      RECT 1.56 1.45 3.59 1.64 ;
      RECT 1.56 0.635 1.75 2.595 ;
      RECT 1.305 2.405 1.75 2.595 ;
  END
END BUFV6_7TV50

MACRO BUFV8_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFV8_7TV50 0 0 ;
  SIZE 10.56 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.525 1.36 1.8 ;
        RECT 0.86 1.525 1.53 1.715 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 2.75 1.355 3.48 ;
        RECT 2.925 2.325 3.205 3.48 ;
        RECT 4.725 2.75 5.005 3.48 ;
        RECT 6.525 2.75 6.805 3.48 ;
        RECT 8.325 2.75 8.605 3.48 ;
        RECT 10.125 2.345 10.405 3.48 ;
        RECT 0 3.24 10.56 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 -0.12 1.405 0.61 ;
        RECT 2.925 -0.12 3.205 0.61 ;
        RECT 4.725 -0.12 5.005 0.565 ;
        RECT 6.525 -0.12 6.805 0.565 ;
        RECT 8.325 -0.12 8.605 0.565 ;
        RECT 10.125 -0.12 10.405 0.61 ;
        RECT 0 -0.12 10.56 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.87 0.595 4.06 0.955 ;
        RECT 5.67 0.595 5.86 0.955 ;
        RECT 6.84 1.52 7.08 1.84 ;
        RECT 6.89 0.765 7.08 2.47 ;
        RECT 7.47 0.595 7.66 0.955 ;
        RECT 9.27 0.595 9.46 0.955 ;
        RECT 3.87 0.765 9.46 0.955 ;
        RECT 3.825 2.28 9.505 2.47 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 10.68 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 11.14 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.27 0.595 0.46 1.015 ;
      RECT 0.27 0.815 2.26 1.015 ;
      RECT 2.07 1.525 6.08 1.715 ;
      RECT 2.07 0.595 2.26 2.47 ;
      RECT 0.225 2.28 2.26 2.47 ;
  END
END BUFV8_7TV50

MACRO BUSHOLD_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUSHOLD_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.815 2.25 2.095 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.915 -0.12 2.195 0.835 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.12 1.52 0.45 1.84 ;
        RECT 0.26 0.595 0.45 2.485 ;
        RECT 0.26 1.805 2.51 1.995 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.54 1.075 3.05 1.265 ;
      RECT 2.86 0.595 3.05 1.27 ;
      RECT 2.71 1.075 2.9 2.485 ;
  END
END BUSHOLD_7TV50

MACRO CLKAND2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 1.065 1.8 ;
        RECT 0.875 1.56 1.065 2.055 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.74 1.56 1.93 2.055 ;
        RECT 1.74 1.56 2.32 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.37 2.315 0.65 3.48 ;
        RECT 1.965 2.97 2.245 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.02 -0.12 2.3 0.83 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.97 0.595 3.16 2.475 ;
        RECT 2.875 2.285 3.16 2.475 ;
        RECT 2.97 1.52 3.24 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.365 0.595 0.555 1.265 ;
      RECT 0.365 1.075 2.675 1.265 ;
      RECT 1.265 1.075 1.455 2.49 ;
  END
END CLKAND2V1_7TV50

MACRO CLKAND2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.38 0.96 3.76 1.34 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.46 1.38 2.76 1.86 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.325 2.4 0.605 3.48 ;
        RECT 2.025 2.4 2.305 3.48 ;
        RECT 3.725 2.4 4.005 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 -0.12 0.505 0.745 ;
        RECT 2.025 -0.12 2.305 0.745 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.56 1.36 1.8 ;
        RECT 1.17 0.51 1.36 2.43 ;
        RECT 1.17 2.24 1.455 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.965 0.555 4.005 0.745 ;
      RECT 1.635 0.99 3.155 1.18 ;
      RECT 2.96 0.99 3.155 2.43 ;
      RECT 2.965 0.555 3.155 2.43 ;
      RECT 2.875 2.24 3.155 2.43 ;
  END
END CLKAND2V2_7TV50

MACRO CLKAND2V3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2V3_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.95 1.84 ;
        RECT 0.76 1.52 0.95 2.04 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.595 1.52 1.785 2.04 ;
        RECT 1.56 1.52 1.845 2.03 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.325 2.4 0.605 3.48 ;
        RECT 2.025 2.4 2.305 3.48 ;
        RECT 3.725 2.79 4.005 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.025 -0.12 2.305 0.83 ;
        RECT 3.825 -0.12 4.105 0.68 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.92 0.64 3.24 0.83 ;
        RECT 3 1.52 3.24 1.84 ;
        RECT 3.05 0.64 3.24 2.44 ;
        RECT 2.875 2.25 4.855 2.44 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.325 0.64 1.36 0.83 ;
      RECT 1.17 1.075 2.68 1.265 ;
      RECT 1.17 0.64 1.36 2.475 ;
      RECT 1.17 2.175 1.41 2.475 ;
  END
END CLKAND2V3_7TV50

MACRO CLKAND2V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2V4_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.515 1.405 0.85 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.505 1.545 1.84 1.975 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 2.4 0.455 3.48 ;
        RECT 1.875 2.4 2.155 3.48 ;
        RECT 3.625 2.79 3.905 3.48 ;
        RECT 5.325 2.4 5.605 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.925 -0.12 2.205 0.73 ;
        RECT 3.725 -0.12 4.005 0.73 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.865 0.595 3.065 1.265 ;
        RECT 4.44 1.075 4.63 2.53 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 2.775 2.34 4.755 2.53 ;
        RECT 4.67 0.595 4.86 1.265 ;
        RECT 2.865 1.075 4.86 1.265 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.225 0.64 1.26 0.83 ;
      RECT 1.07 1.155 2.595 1.345 ;
      RECT 1.07 0.64 1.26 2.59 ;
  END
END CLKAND2V4_7TV50

MACRO CLKBUFV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFV1_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.875 1.56 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.545 1.345 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 -0.12 1.345 0.875 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.01 0.595 2.2 2.475 ;
        RECT 2.01 1.52 2.28 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.21 1.805 1.72 1.995 ;
      RECT 0.21 0.595 0.4 2.475 ;
  END
END CLKBUFV1_7TV50

MACRO CLKBUFV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFV2_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.75 1.04 1.32 1.36 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 2.195 1.405 3.48 ;
        RECT 2.84 2.36 3.12 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 -0.12 1.405 0.83 ;
        RECT 2.925 -0.12 3.205 0.83 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.07 0.595 2.26 2.475 ;
        RECT 1.99 2.195 2.26 2.475 ;
        RECT 2.04 1.52 2.28 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.27 0.595 0.46 1.995 ;
      RECT 0.27 1.805 1.78 1.995 ;
      RECT 0.32 1.805 0.51 2.475 ;
  END
END CLKBUFV2_7TV50

MACRO CLKBUFV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFV3_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.9 1.52 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 2.36 1.335 3.48 ;
        RECT 2.85 2.795 3.13 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 2.855 -0.12 3.135 0.81 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.595 2.19 2.43 ;
        RECT 2 1.52 2.28 1.84 ;
        RECT 2 2.24 3.98 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.805 1.71 1.995 ;
      RECT 0.2 0.595 0.39 2.475 ;
  END
END CLKBUFV3_7TV50

MACRO CLKBUFV4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFV4_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.84 2.12 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.565 0.435 3.48 ;
        RECT 1.925 2.565 2.205 3.48 ;
        RECT 3.625 2.75 3.905 3.48 ;
        RECT 5.325 2.36 5.605 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.925 -0.12 2.205 0.875 ;
        RECT 3.725 -0.12 4.005 0.83 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.87 0.595 3.06 1.225 ;
        RECT 4.44 1.52 4.755 1.84 ;
        RECT 4.565 1.035 4.755 2.43 ;
        RECT 2.775 2.24 4.755 2.43 ;
        RECT 4.67 0.595 4.86 1.225 ;
        RECT 2.87 1.035 4.86 1.225 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.025 0.64 1.31 0.83 ;
      RECT 1.12 1.805 3.525 1.995 ;
      RECT 1.12 0.64 1.31 2.475 ;
  END
END CLKBUFV4_7TV50

MACRO CLKBUFV6_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFV6_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.975 1.84 ;
        RECT 0.7 1.52 0.975 2.04 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.325 2.29 0.605 3.48 ;
        RECT 2.025 2.29 2.305 3.48 ;
        RECT 3.725 2.745 4.005 3.48 ;
        RECT 5.425 2.745 5.705 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 -0.12 0.505 0.875 ;
        RECT 2.025 -0.12 2.305 0.875 ;
        RECT 3.825 -0.12 4.105 0.835 ;
        RECT 5.625 -0.12 5.905 0.875 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.97 0.595 3.16 1.225 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.49 1.035 4.68 2.51 ;
        RECT 4.77 0.595 4.96 1.225 ;
        RECT 2.97 1.035 4.96 1.225 ;
        RECT 2.875 2.32 6.555 2.51 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.17 0.595 1.36 1.04 ;
      RECT 1.22 0.84 1.425 1.615 ;
      RECT 1.22 1.425 3.64 1.615 ;
      RECT 1.22 0.84 1.415 2.635 ;
  END
END CLKBUFV6_7TV50

MACRO CLKBUFV8_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFV8_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.53 1.04 0.84 1.61 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.75 1.285 3.48 ;
        RECT 2.705 2.36 2.985 3.48 ;
        RECT 4.405 2.795 4.685 3.48 ;
        RECT 6.105 2.795 6.385 3.48 ;
        RECT 7.805 2.795 8.085 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.905 -0.12 1.185 0.83 ;
        RECT 2.705 -0.12 2.985 0.875 ;
        RECT 4.565 -0.12 4.845 0.44 ;
        RECT 6.425 -0.12 6.705 0.875 ;
        RECT 8.225 -0.12 8.505 0.83 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.605 0.64 5.805 0.83 ;
        RECT 5.615 0.64 5.805 2.455 ;
        RECT 7.32 1.52 7.56 1.84 ;
        RECT 7.37 0.595 7.56 2.455 ;
        RECT 3.555 2.265 8.935 2.455 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.85 0.595 2.04 2.495 ;
      RECT 1.85 1.67 5.11 1.86 ;
      RECT 1.85 1.67 2.045 2.495 ;
      RECT 0.155 2.295 2.135 2.495 ;
  END
END CLKBUFV8_7TV50

MACRO CLKINV16_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV16_7TV50 0 0 ;
  SIZE 12.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.97 ;
        RECT 4.18 1.78 5.24 1.97 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.405 0.565 3.48 ;
        RECT 1.985 2.795 2.265 3.48 ;
        RECT 3.685 2.795 3.965 3.48 ;
        RECT 5.385 2.795 5.665 3.48 ;
        RECT 7.085 2.795 7.365 3.48 ;
        RECT 8.785 2.795 9.065 3.48 ;
        RECT 10.485 2.795 10.765 3.48 ;
        RECT 12.185 2.405 12.465 3.48 ;
        RECT 0 3.24 12.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.185 -0.12 1.465 0.83 ;
        RECT 2.985 -0.12 3.265 0.83 ;
        RECT 4.785 -0.12 5.065 0.83 ;
        RECT 6.585 -0.12 6.865 0.83 ;
        RECT 8.385 -0.12 8.665 0.83 ;
        RECT 10.185 -0.12 10.465 0.83 ;
        RECT 11.985 -0.12 12.265 0.83 ;
        RECT 0 -0.12 12.96 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.595 0.52 1.22 ;
        RECT 2.13 0.595 2.32 1.22 ;
        RECT 3.93 0.595 4.12 1.22 ;
        RECT 5.73 0.595 5.92 1.22 ;
        RECT 6.28 1.03 6.47 2.5 ;
        RECT 6.28 1.52 6.6 1.84 ;
        RECT 7.53 0.595 7.72 1.22 ;
        RECT 9.33 0.595 9.52 1.22 ;
        RECT 11.13 0.595 11.32 1.22 ;
        RECT 0.33 1.03 11.32 1.22 ;
        RECT 1.135 2.31 11.615 2.5 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 13.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 13.54 3.94 ;
    END
  END VNW
END CLKINV16_7TV50

MACRO CLKINV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV1_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.52 1.52 0.84 1.97 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.36 0.435 3.48 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.83 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.05 1.04 1.24 2.475 ;
        RECT 1.1 0.55 1.29 1.36 ;
        RECT 1.05 1.04 1.32 1.36 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
END CLKINV1_7TV50

MACRO CLKINV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV2_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.04 0.84 1.36 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.36 0.485 3.48 ;
        RECT 1.905 2.36 2.185 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.84 ;
        RECT 1.955 -0.12 2.235 0.84 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.56 1.29 2.64 ;
        RECT 1.08 1.04 1.32 1.36 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
END CLKINV2_7TV50

MACRO CLKINV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV3_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.885 1.52 1.32 1.94 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.36 2.36 0.64 3.48 ;
        RECT 2.06 2.75 2.34 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.36 -0.12 0.64 0.81 ;
        RECT 2.16 -0.12 2.44 0.81 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.305 0.595 1.495 1.285 ;
        RECT 1.305 1.095 1.81 1.285 ;
        RECT 1.56 1.52 1.81 1.84 ;
        RECT 1.62 1.095 1.81 2.55 ;
        RECT 1.62 2.355 3.19 2.55 ;
        RECT 1.21 2.36 3.19 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
END CLKINV3_7TV50

MACRO CLKINV4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV4_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.84 2.04 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.455 2.36 0.735 3.48 ;
        RECT 2.155 2.795 2.435 3.48 ;
        RECT 3.855 2.36 4.135 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.555 -0.12 1.845 0.83 ;
        RECT 3.365 -0.12 3.645 0.865 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.71 0.595 0.9 1.22 ;
        RECT 0.71 1.03 2.7 1.22 ;
        RECT 2.51 0.595 2.7 2.43 ;
        RECT 2.51 1.52 2.76 1.84 ;
        RECT 1.305 2.24 3.49 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
END CLKINV4_7TV50

MACRO CLKINV6_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV6_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.52 2.28 1.84 ;
        RECT 1.445 1.65 2.51 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.36 0.435 3.48 ;
        RECT 1.855 2.75 2.135 3.48 ;
        RECT 3.555 2.75 3.835 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.555 -0.12 0.835 0.82 ;
        RECT 2.355 -0.12 2.635 0.775 ;
        RECT 4.155 -0.12 4.435 0.82 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5 0.59 1.69 1.165 ;
        RECT 3 0.975 3.19 2.43 ;
        RECT 3 1.52 3.24 1.84 ;
        RECT 3.3 0.59 3.49 1.165 ;
        RECT 1.5 0.975 3.49 1.165 ;
        RECT 1.005 2.24 4.705 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
END CLKINV6_7TV50

MACRO CLKINV8_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINV8_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.8 1.84 ;
        RECT 1.525 1.56 2.605 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.1 2.745 1.38 3.48 ;
        RECT 2.8 2.745 3.08 3.48 ;
        RECT 4.5 2.745 4.78 3.48 ;
        RECT 6.2 2.7 6.48 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.25 -0.12 0.53 0.855 ;
        RECT 2.05 -0.12 2.33 0.81 ;
        RECT 3.85 -0.12 4.13 0.81 ;
        RECT 5.65 -0.12 5.93 0.855 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.195 0.595 1.385 1.2 ;
        RECT 2.995 0.595 3.185 1.2 ;
        RECT 3 1.01 3.19 2.48 ;
        RECT 3 1.52 3.24 1.84 ;
        RECT 4.795 0.595 4.985 1.2 ;
        RECT 1.195 1.01 4.985 1.2 ;
        RECT 0.25 2.29 5.63 2.48 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
END CLKINV8_7TV50

MACRO CLKLAHAQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLAHAQV1_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.225 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.56 3.24 1.225 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.6 0.6 12.28 0.84 ;
        RECT 12.09 0.6 12.28 2.48 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.88 1.56 8.56 1.8 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.25 1.285 3.48 ;
        RECT 2.445 2.235 2.725 3.48 ;
        RECT 5.705 2.97 5.985 3.48 ;
        RECT 8.1 2.55 8.335 3.48 ;
        RECT 11.195 2.795 11.475 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.79 ;
        RECT 2.545 -0.12 2.78 0.79 ;
        RECT 5.945 -0.12 6.225 0.79 ;
        RECT 8.335 -0.12 8.615 0.935 ;
        RECT 10.995 -0.12 11.275 0.83 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.075 1.46 ;
        RECT -0.12 -0.24 12.6 1.375 ;
        RECT 6.98 -0.24 10.575 1.565 ;
        RECT 6.98 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.075 1.375 6.98 3.94 ;
        RECT -0.58 1.46 6.98 3.94 ;
        RECT 10.575 1.46 13.06 3.94 ;
        RECT -0.58 1.565 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.645 1.66 1.835 ;
      RECT 0.2 0.51 0.39 2.475 ;
      RECT 4.29 1.675 6.42 1.865 ;
      RECT 4.29 0.51 4.48 2.535 ;
      RECT 4.045 2.345 4.48 2.535 ;
      RECT 6.89 0.51 7.08 1.18 ;
      RECT 5.57 0.99 7.08 1.18 ;
      RECT 6.705 0.99 6.895 2.535 ;
      RECT 6.615 2.345 6.895 2.535 ;
      RECT 7.48 0.7 7.67 1.325 ;
      RECT 7.295 1.135 8.945 1.325 ;
      RECT 8.755 1.135 8.945 1.415 ;
      RECT 7.295 1.135 7.485 2.535 ;
      RECT 7.205 2.345 7.485 2.535 ;
      RECT 3.44 0.99 4 1.18 ;
      RECT 2 1.63 3.63 1.82 ;
      RECT 8.855 1.99 10.25 2.18 ;
      RECT 7.71 2.16 9.045 2.35 ;
      RECT 2 0.51 2.19 2.43 ;
      RECT 1.855 2.24 2.19 2.43 ;
      RECT 4.885 2.58 6.415 2.77 ;
      RECT 6.225 2.58 6.415 2.965 ;
      RECT 3.44 0.99 3.63 2.98 ;
      RECT 7.71 2.16 7.9 2.965 ;
      RECT 6.225 2.775 7.9 2.965 ;
      RECT 4.885 2.58 5.075 2.98 ;
      RECT 3.44 2.79 5.075 2.98 ;
      RECT 8.95 2.67 9.14 3.005 ;
      RECT 10.345 2.795 10.625 3.005 ;
      RECT 8.95 2.815 10.625 3.005 ;
      RECT 9.705 1.135 9.895 1.655 ;
      RECT 9.705 1.465 10.955 1.655 ;
      RECT 10.765 1.465 10.955 2.18 ;
      RECT 10.14 0.595 10.33 1.265 ;
      RECT 10.14 1.075 11.65 1.265 ;
      RECT 11.155 1.075 11.345 2.57 ;
      RECT 9.495 2.38 11.345 2.57 ;
      RECT 9.495 2.38 9.775 2.615 ;
  END
END CLKLAHAQV1_7TV50

MACRO CLKLAHAQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLAHAQV2_7TV50 0 0 ;
  SIZE 15.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.205 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.56 3.24 1.16 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.18 0.585 14.24 0.84 ;
        RECT 14.05 0.585 14.24 2.475 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.76 1.56 8.36 1.8 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.21 1.285 3.48 ;
        RECT 2.445 2.195 2.725 3.48 ;
        RECT 5.705 2.655 5.985 3.48 ;
        RECT 8.1 2.535 8.335 3.48 ;
        RECT 9.755 2.79 10.035 3.48 ;
        RECT 13.155 2.275 13.435 3.48 ;
        RECT 14.855 2.275 15.135 3.48 ;
        RECT 0 3.24 15.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.69 ;
        RECT 2.545 -0.12 2.78 0.655 ;
        RECT 5.945 -0.12 6.225 0.69 ;
        RECT 7.775 -0.12 8.055 0.565 ;
        RECT 9.605 -0.12 9.885 0.565 ;
        RECT 12.325 -0.12 12.56 0.61 ;
        RECT 0 -0.12 15.36 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.935 1.46 ;
        RECT -0.12 -0.24 15.48 1.275 ;
        RECT 6.405 -0.24 9.32 1.53 ;
        RECT 6.405 -0.24 15.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 1.935 1.275 6.405 3.94 ;
        RECT -0.58 1.46 6.405 3.94 ;
        RECT 9.32 1.46 15.94 3.94 ;
        RECT -0.58 1.53 15.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.645 1.66 1.835 ;
      RECT 0.2 0.49 0.39 2.475 ;
      RECT 6.905 0.71 7.185 0.9 ;
      RECT 6.905 0.71 7.095 1.83 ;
      RECT 5.27 1.64 7.095 1.83 ;
      RECT 6.705 1.64 6.895 2.5 ;
      RECT 6.615 2.31 6.895 2.5 ;
      RECT 8.735 0.71 9.015 0.9 ;
      RECT 8.825 0.71 9.015 1.36 ;
      RECT 7.295 1.17 9.56 1.36 ;
      RECT 7.295 1.17 7.485 2.52 ;
      RECT 7.205 2.33 7.485 2.52 ;
      RECT 6.465 0.32 7.575 0.51 ;
      RECT 8.255 0.32 9.405 0.51 ;
      RECT 7.385 0.32 7.575 0.955 ;
      RECT 9.215 0.32 9.405 0.955 ;
      RECT 8.255 0.32 8.445 0.955 ;
      RECT 7.385 0.765 8.445 0.955 ;
      RECT 9.215 0.765 11.015 0.955 ;
      RECT 10.825 0.765 11.015 1.045 ;
      RECT 6.465 0.32 6.655 1.08 ;
      RECT 4.29 0.89 6.655 1.08 ;
      RECT 4.29 0.41 4.48 2.5 ;
      RECT 4.045 2.31 4.48 2.5 ;
      RECT 3.44 0.89 4 1.08 ;
      RECT 2 0.41 2.19 1.76 ;
      RECT 1.9 1.57 3.63 1.76 ;
      RECT 8.56 1.895 11.735 2.085 ;
      RECT 11.545 0.765 11.735 2.085 ;
      RECT 7.71 2.075 8.75 2.265 ;
      RECT 4.885 2.265 6.415 2.455 ;
      RECT 1.9 1.57 2.09 2.475 ;
      RECT 6.225 2.265 6.415 2.92 ;
      RECT 3.44 0.89 3.63 2.945 ;
      RECT 7.71 2.075 7.9 2.92 ;
      RECT 6.225 2.73 7.9 2.92 ;
      RECT 4.885 2.265 5.075 2.945 ;
      RECT 3.44 2.755 5.075 2.945 ;
      RECT 8.905 2.4 10.84 2.59 ;
      RECT 10.65 2.4 10.84 2.91 ;
      RECT 10.65 2.72 12.585 2.91 ;
      RECT 11.365 0.375 12.125 0.565 ;
      RECT 11.935 1.805 13.81 1.995 ;
      RECT 11.935 0.375 12.125 2.52 ;
      RECT 11.455 2.33 12.125 2.52 ;
  END
END CLKLAHAQV2_7TV50

MACRO CLKLAHAQV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLAHAQV3_7TV50 0 0 ;
  SIZE 16.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.16 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.56 3.24 1.16 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.05 1.965 14.24 2.475 ;
        RECT 14.95 0.51 15.14 2.155 ;
        RECT 14.95 0.51 15.24 0.88 ;
        RECT 14.05 1.965 15.94 2.155 ;
        RECT 15.75 1.965 15.94 2.475 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.76 1.56 8.36 1.8 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.32 1.285 3.48 ;
        RECT 2.445 2.195 2.725 3.48 ;
        RECT 5.705 2.655 5.985 3.48 ;
        RECT 8.1 2.535 8.335 3.48 ;
        RECT 9.755 2.79 10.035 3.48 ;
        RECT 13.155 2.275 13.435 3.48 ;
        RECT 14.855 2.355 15.135 3.48 ;
        RECT 0 3.24 16.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.69 ;
        RECT 2.545 -0.12 2.78 0.655 ;
        RECT 5.945 -0.12 6.225 0.69 ;
        RECT 7.775 -0.12 8.055 0.565 ;
        RECT 9.605 -0.12 9.885 0.565 ;
        RECT 12.325 -0.12 12.56 0.61 ;
        RECT 14.005 -0.12 14.285 0.79 ;
        RECT 15.805 -0.12 16.085 0.745 ;
        RECT 0 -0.12 16.32 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.935 1.46 ;
        RECT -0.12 -0.24 16.44 1.275 ;
        RECT 6.405 -0.24 9.32 1.53 ;
        RECT 6.405 -0.24 16.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 1.935 1.275 6.405 3.94 ;
        RECT -0.58 1.46 6.405 3.94 ;
        RECT 9.32 1.46 16.9 3.94 ;
        RECT -0.58 1.53 16.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.645 1.66 1.835 ;
      RECT 0.2 0.41 0.39 2.475 ;
      RECT 6.905 0.71 7.185 0.9 ;
      RECT 6.905 0.71 7.095 1.83 ;
      RECT 5.27 1.64 7.095 1.83 ;
      RECT 6.705 1.64 6.895 2.5 ;
      RECT 6.615 2.31 6.895 2.5 ;
      RECT 8.735 0.71 9.015 0.9 ;
      RECT 8.825 0.71 9.015 1.36 ;
      RECT 7.295 1.17 9.56 1.36 ;
      RECT 7.295 1.17 7.485 2.52 ;
      RECT 7.205 2.33 7.485 2.52 ;
      RECT 6.465 0.32 7.575 0.51 ;
      RECT 8.255 0.32 9.405 0.51 ;
      RECT 7.385 0.32 7.575 0.955 ;
      RECT 9.215 0.32 9.405 0.955 ;
      RECT 8.255 0.32 8.445 0.955 ;
      RECT 7.385 0.765 8.445 0.955 ;
      RECT 9.215 0.765 11.015 0.955 ;
      RECT 10.825 0.765 11.015 1.045 ;
      RECT 6.465 0.32 6.655 1.08 ;
      RECT 4.29 0.89 6.655 1.08 ;
      RECT 4.29 0.41 4.48 2.5 ;
      RECT 4.045 2.31 4.48 2.5 ;
      RECT 3.44 0.89 4 1.08 ;
      RECT 2 0.41 2.19 1.82 ;
      RECT 1.9 1.63 3.63 1.82 ;
      RECT 8.56 1.895 11.735 2.085 ;
      RECT 11.545 0.765 11.735 2.085 ;
      RECT 7.71 2.075 8.75 2.265 ;
      RECT 4.885 2.265 6.415 2.455 ;
      RECT 1.9 1.63 2.09 2.475 ;
      RECT 6.225 2.265 6.415 2.92 ;
      RECT 3.44 0.89 3.63 2.945 ;
      RECT 7.71 2.075 7.9 2.92 ;
      RECT 6.225 2.73 7.9 2.92 ;
      RECT 4.885 2.265 5.075 2.945 ;
      RECT 3.44 2.755 5.075 2.945 ;
      RECT 8.905 2.4 10.84 2.59 ;
      RECT 10.65 2.4 10.84 2.91 ;
      RECT 10.65 2.72 12.585 2.91 ;
      RECT 11.365 0.375 12.125 0.565 ;
      RECT 11.935 1.575 14.46 1.765 ;
      RECT 11.935 0.375 12.125 2.52 ;
      RECT 11.455 2.33 12.125 2.52 ;
  END
END CLKLAHAQV3_7TV50

MACRO CLKLAHQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLAHQV1_7TV50 0 0 ;
  SIZE 12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 1.05 1.36 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.85 1 4.245 1.37 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.12 0.6 11.66 0.84 ;
        RECT 11.47 0.6 11.66 2.48 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.895 1 3.345 1.37 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.25 1.285 3.48 ;
        RECT 2.765 2.405 3.045 3.48 ;
        RECT 6.81 2.97 7.09 3.48 ;
        RECT 10.575 2.795 10.855 3.48 ;
        RECT 0 3.24 12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.79 ;
        RECT 3.49 -0.12 3.77 0.79 ;
        RECT 7.025 -0.12 7.305 0.79 ;
        RECT 8.515 -0.12 8.795 0.935 ;
        RECT 10.375 -0.12 10.655 0.83 ;
        RECT 0 -0.12 12 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.075 1.46 ;
        RECT -0.12 -0.24 12.12 1.375 ;
        RECT 8.06 -0.24 9.955 1.565 ;
        RECT 8.06 -0.24 12.12 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.075 1.375 8.06 3.94 ;
        RECT -0.58 1.46 8.06 3.94 ;
        RECT 9.955 1.46 12.58 3.94 ;
        RECT -0.58 1.565 12.58 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.805 1.66 1.995 ;
      RECT 0.2 0.51 0.39 2.475 ;
      RECT 2.505 0.555 2.825 0.745 ;
      RECT 2.505 0.555 2.695 1.76 ;
      RECT 4.445 0.505 4.635 1.76 ;
      RECT 2.505 1.57 4.635 1.76 ;
      RECT 5.37 1.95 7.525 2.14 ;
      RECT 5.37 0.51 5.56 2.585 ;
      RECT 5.15 2.395 5.56 2.585 ;
      RECT 7.97 0.51 8.16 1.18 ;
      RECT 6.635 0.99 8.16 1.18 ;
      RECT 7.81 0.99 8 2.575 ;
      RECT 7.72 2.385 8 2.575 ;
      RECT 4.845 0.945 5.035 2.205 ;
      RECT 2 2.015 5.035 2.205 ;
      RECT 2 0.51 2.19 2.43 ;
      RECT 1.855 2.24 2.19 2.43 ;
      RECT 8.26 2.35 9.53 2.54 ;
      RECT 5.99 2.58 7.52 2.77 ;
      RECT 7.33 2.58 7.52 2.965 ;
      RECT 4.52 2.015 4.71 3.03 ;
      RECT 8.26 2.35 8.45 2.965 ;
      RECT 7.33 2.775 8.45 2.965 ;
      RECT 5.99 2.58 6.18 3.03 ;
      RECT 4.52 2.84 6.18 3.03 ;
      RECT 9.085 1.135 9.275 1.655 ;
      RECT 9.085 1.465 10.335 1.655 ;
      RECT 10.145 1.465 10.335 2.18 ;
      RECT 9.52 0.595 9.71 1.265 ;
      RECT 9.52 1.075 11.03 1.265 ;
      RECT 10.535 1.075 10.725 2.57 ;
      RECT 10.01 2.38 10.725 2.57 ;
      RECT 10.01 2.38 10.2 2.975 ;
      RECT 8.875 2.785 10.2 2.975 ;
  END
END CLKLAHQV1_7TV50

MACRO CLKLAHQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLAHQV2_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 1.05 1.36 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.85 1 4.245 1.37 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.095 1.56 11.285 2.48 ;
        RECT 11.315 0.595 11.505 1.8 ;
        RECT 11.095 1.56 11.505 1.8 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.895 1 3.345 1.37 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.25 1.285 3.48 ;
        RECT 2.765 2.405 3.045 3.48 ;
        RECT 6.81 2.97 7.09 3.48 ;
        RECT 10.2 2.795 10.48 3.48 ;
        RECT 11.9 2.405 12.185 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.79 ;
        RECT 3.49 -0.12 3.77 0.79 ;
        RECT 7.025 -0.12 7.305 0.79 ;
        RECT 8.515 -0.12 8.795 0.745 ;
        RECT 10.37 -0.12 10.65 0.745 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.075 1.46 ;
        RECT -0.12 -0.24 12.6 1.375 ;
        RECT 8.06 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.075 1.375 8.06 3.94 ;
        RECT -0.58 1.46 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.805 1.66 1.995 ;
      RECT 0.2 0.51 0.39 2.475 ;
      RECT 2.505 0.555 2.825 0.745 ;
      RECT 2.505 0.555 2.695 1.76 ;
      RECT 4.445 0.505 4.635 1.76 ;
      RECT 2.505 1.57 4.635 1.76 ;
      RECT 5.37 1.95 7.525 2.14 ;
      RECT 5.37 0.51 5.56 2.585 ;
      RECT 5.15 2.395 5.56 2.585 ;
      RECT 7.97 0.51 8.16 1.18 ;
      RECT 6.635 0.99 8.16 1.18 ;
      RECT 7.765 0.99 7.955 2.62 ;
      RECT 8.155 1.81 9.155 2 ;
      RECT 4.845 0.945 5.035 2.205 ;
      RECT 2 2.015 5.035 2.205 ;
      RECT 2 0.51 2.19 2.43 ;
      RECT 1.855 2.24 2.19 2.43 ;
      RECT 5.99 2.58 7.52 2.77 ;
      RECT 7.33 2.58 7.52 3.01 ;
      RECT 4.52 2.015 4.71 3.03 ;
      RECT 8.155 1.81 8.345 3.01 ;
      RECT 7.33 2.82 8.345 3.01 ;
      RECT 5.99 2.58 6.18 3.03 ;
      RECT 4.52 2.84 6.18 3.03 ;
      RECT 9.085 0.925 9.275 1.57 ;
      RECT 9.085 1.38 9.655 1.57 ;
      RECT 9.465 1.52 10.315 1.71 ;
      RECT 9.47 0.555 10.17 0.745 ;
      RECT 9.98 0.555 10.17 1.265 ;
      RECT 9.98 1.075 11.08 1.265 ;
      RECT 8.545 2.205 8.74 2.44 ;
      RECT 10.595 1.075 10.785 2.44 ;
      RECT 8.545 2.245 10.785 2.44 ;
      RECT 8.545 2.205 8.735 2.485 ;
  END
END CLKLAHQV2_7TV50

MACRO CLKLAHQV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLAHQV3_7TV50 0 0 ;
  SIZE 12.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 1.05 1.36 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.85 1 4.245 1.37 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.81 1.56 11 2.48 ;
        RECT 11.57 0.595 11.76 1.8 ;
        RECT 10.81 1.56 11.76 1.8 ;
        RECT 10.81 1.61 12.7 1.8 ;
        RECT 12.51 1.61 12.7 2.48 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.895 1 3.345 1.37 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.25 1.285 3.48 ;
        RECT 2.505 2.405 2.785 3.48 ;
        RECT 6.525 2.97 6.805 3.48 ;
        RECT 9.915 2.795 10.195 3.48 ;
        RECT 11.615 2.405 11.9 3.48 ;
        RECT 0 3.24 12.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.79 ;
        RECT 3.49 -0.12 3.77 0.79 ;
        RECT 7.025 -0.12 7.305 0.79 ;
        RECT 8.515 -0.12 8.795 0.745 ;
        RECT 10.67 -0.12 10.86 0.79 ;
        RECT 12.425 -0.12 12.705 0.745 ;
        RECT 0 -0.12 12.96 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.075 1.46 ;
        RECT -0.12 -0.24 13.08 1.375 ;
        RECT 7.775 -0.24 13.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.075 1.375 7.775 3.94 ;
        RECT -0.58 1.46 13.54 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.805 1.66 1.995 ;
      RECT 0.2 0.51 0.39 2.475 ;
      RECT 2.505 0.555 2.825 0.745 ;
      RECT 2.505 0.555 2.695 1.76 ;
      RECT 4.445 0.505 4.635 1.76 ;
      RECT 2.505 1.57 4.635 1.76 ;
      RECT 5.37 1.95 7.24 2.14 ;
      RECT 5.37 0.51 5.56 2.585 ;
      RECT 4.835 2.395 5.56 2.585 ;
      RECT 7.97 0.51 8.16 1.18 ;
      RECT 6.635 0.99 8.16 1.18 ;
      RECT 7.48 0.99 7.67 2.62 ;
      RECT 9.89 0.945 10.08 2 ;
      RECT 7.87 1.81 10.08 2 ;
      RECT 4.845 0.945 5.035 2.185 ;
      RECT 2 1.995 5.035 2.185 ;
      RECT 2 0.51 2.19 2.43 ;
      RECT 1.855 2.22 2.19 2.43 ;
      RECT 5.765 2.58 7.235 2.77 ;
      RECT 7.045 2.58 7.235 3.01 ;
      RECT 4.26 1.995 4.45 3.03 ;
      RECT 7.87 1.81 8.06 3.01 ;
      RECT 7.045 2.82 8.06 3.01 ;
      RECT 5.765 2.58 5.955 3.03 ;
      RECT 4.26 2.84 5.955 3.03 ;
      RECT 9.46 0.555 10.47 0.745 ;
      RECT 10.28 1.075 11.335 1.265 ;
      RECT 10.28 0.555 10.47 2.44 ;
      RECT 8.36 2.245 10.47 2.44 ;
      RECT 8.36 2.205 8.55 2.485 ;
  END
END CLKLAHQV3_7TV50

MACRO CLKLANAQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLANAQV1_7TV50 0 0 ;
  SIZE 13.44 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.345 1.51 1.8 1.85 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.455 3.325 1.9 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.165 2.04 12.355 2.48 ;
        RECT 12.775 0.52 12.965 2.28 ;
        RECT 12.165 2.04 12.965 2.28 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.68 1.04 11.16 1.425 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.97 1.345 3.48 ;
        RECT 2.655 2.97 2.935 3.48 ;
        RECT 6.865 2.355 7.125 3.48 ;
        RECT 8.71 2.795 8.99 3.48 ;
        RECT 11.255 2.79 11.535 3.48 ;
        RECT 0 3.24 13.44 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 -0.12 1.355 0.565 ;
        RECT 3.465 -0.12 3.745 0.64 ;
        RECT 3.465 -0.12 7.145 0.195 ;
        RECT 6.865 -0.12 7.145 0.64 ;
        RECT 10.34 -0.12 10.62 0.39 ;
        RECT 11.83 -0.12 12.11 0.76 ;
        RECT 0 -0.12 13.44 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.095 1.46 ;
        RECT -0.12 -0.24 13.56 1.27 ;
        RECT 3.3 -0.24 13.56 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 1.095 1.27 3.3 3.94 ;
        RECT -0.58 1.46 14.02 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.065 0.885 4.97 1.075 ;
      RECT 0.675 1.96 0.865 2.38 ;
      RECT 2.065 0.33 2.255 2.38 ;
      RECT 0.675 2.19 2.315 2.38 ;
      RECT 5.21 0.935 7.52 1.125 ;
      RECT 5.21 0.405 5.4 2.445 ;
      RECT 4.315 2.255 5.4 2.445 ;
      RECT 5.68 1.9 7.515 2.09 ;
      RECT 8.24 1.9 9.165 2.09 ;
      RECT 0.2 0.33 0.39 2.77 ;
      RECT 3.925 1.76 4.115 2.835 ;
      RECT 7.325 1.9 7.515 2.93 ;
      RECT 0.2 2.58 4.115 2.77 ;
      RECT 5.68 1.35 5.87 2.835 ;
      RECT 3.925 2.645 5.87 2.835 ;
      RECT 8.24 1.9 8.43 2.93 ;
      RECT 7.325 2.74 8.43 2.93 ;
      RECT 7.81 0.4 8 1.7 ;
      RECT 6.43 1.51 10.04 1.7 ;
      RECT 7.805 1.51 7.995 2.435 ;
      RECT 7.715 2.24 7.995 2.435 ;
      RECT 9.425 0.39 9.615 0.795 ;
      RECT 10.975 0.515 11.165 0.795 ;
      RECT 9.425 0.605 11.165 0.795 ;
      RECT 8.525 0.52 8.715 1.31 ;
      RECT 8.525 1.12 10.43 1.31 ;
      RECT 10.24 1.12 10.43 2.205 ;
      RECT 11.69 1.765 11.88 2.205 ;
      RECT 9.61 2.015 11.88 2.205 ;
      RECT 9.61 2.015 9.8 3.01 ;
  END
END CLKLANAQV1_7TV50

MACRO CLKLANAQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLANAQV2_7TV50 0 0 ;
  SIZE 13.44 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.345 1.51 1.8 1.85 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.455 3.325 1.9 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.175 2.04 12.365 2.61 ;
        RECT 12.845 0.35 13.035 2.28 ;
        RECT 12.175 2.04 13.035 2.28 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.68 1.04 11.16 1.425 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.97 1.345 3.48 ;
        RECT 2.655 2.97 2.935 3.48 ;
        RECT 6.865 2.54 7.125 3.48 ;
        RECT 8.71 2.795 8.99 3.48 ;
        RECT 11.255 2.79 11.535 3.48 ;
        RECT 12.98 2.795 13.26 3.48 ;
        RECT 0 3.24 13.44 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 -0.12 1.355 0.565 ;
        RECT 3.465 -0.12 3.745 0.565 ;
        RECT 6.865 -0.12 7.145 0.565 ;
        RECT 10.34 -0.12 10.62 0.39 ;
        RECT 11.89 -0.12 12.19 0.57 ;
        RECT 0 -0.12 13.44 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.095 1.46 ;
        RECT -0.12 -0.24 13.56 1.27 ;
        RECT 3.3 -0.24 13.56 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 1.095 1.27 3.3 3.94 ;
        RECT -0.58 1.46 14.02 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.065 0.81 4.97 1 ;
      RECT 0.675 1.96 0.865 2.38 ;
      RECT 2.065 0.33 2.255 2.38 ;
      RECT 0.675 2.19 2.315 2.38 ;
      RECT 5.21 0.86 7.52 1.05 ;
      RECT 5.21 0.33 5.4 2.63 ;
      RECT 4.315 2.44 5.4 2.63 ;
      RECT 8.24 1.9 9.165 2.09 ;
      RECT 5.735 2.085 7.515 2.275 ;
      RECT 0.2 0.33 0.39 2.77 ;
      RECT 0.2 2.58 4.075 2.77 ;
      RECT 3.885 1.945 4.075 3.02 ;
      RECT 7.325 2.085 7.515 3.04 ;
      RECT 5.735 1.275 5.925 3.02 ;
      RECT 3.885 2.83 5.925 3.02 ;
      RECT 8.24 1.9 8.43 3.04 ;
      RECT 7.325 2.85 8.43 3.04 ;
      RECT 7.81 0.325 8 1.7 ;
      RECT 7.81 1.51 10.02 1.7 ;
      RECT 6.43 1.64 7.995 1.83 ;
      RECT 7.805 1.64 7.995 2.62 ;
      RECT 7.715 2.425 7.995 2.62 ;
      RECT 9.425 0.35 9.615 0.795 ;
      RECT 11.045 0.39 11.235 0.795 ;
      RECT 9.425 0.605 11.235 0.795 ;
      RECT 8.525 0.39 8.715 1.31 ;
      RECT 8.525 1.12 10.43 1.31 ;
      RECT 10.24 1.12 10.43 2.205 ;
      RECT 11.785 1.765 11.975 2.205 ;
      RECT 9.61 2.015 11.975 2.205 ;
      RECT 9.61 2.015 9.8 2.66 ;
  END
END CLKLANAQV2_7TV50

MACRO CLKLANAQV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLANAQV3_7TV50 0 0 ;
  SIZE 14.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.345 1.51 1.84 1.85 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.455 3.325 1.9 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.8 0.395 13.5 0.585 ;
        RECT 13.31 0.395 13.5 2.435 ;
        RECT 13.31 2 13.8 2.435 ;
        RECT 12.13 2.245 14.11 2.435 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.68 1.04 11.16 1.425 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.97 1.345 3.48 ;
        RECT 2.655 2.97 2.935 3.48 ;
        RECT 6.865 2.52 7.125 3.48 ;
        RECT 8.71 2.355 8.99 3.48 ;
        RECT 11.255 2.405 11.535 3.48 ;
        RECT 12.98 2.795 13.26 3.48 ;
        RECT 0 3.24 14.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.12 -0.12 1.31 0.61 ;
        RECT 3.465 -0.12 3.745 0.565 ;
        RECT 6.865 -0.12 7.145 0.565 ;
        RECT 10.34 -0.12 10.62 0.39 ;
        RECT 11.9 -0.12 12.18 0.565 ;
        RECT 13.7 -0.12 13.98 0.565 ;
        RECT 0 -0.12 14.4 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.095 1.46 ;
        RECT -0.12 -0.24 14.52 1.27 ;
        RECT 3.3 -0.24 14.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 1.095 1.27 3.3 3.94 ;
        RECT -0.58 1.46 14.98 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.065 0.86 4.97 1.05 ;
      RECT 0.59 1.96 0.78 2.38 ;
      RECT 2.065 0.33 2.255 2.38 ;
      RECT 0.59 2.19 2.315 2.38 ;
      RECT 5.21 0.81 7.525 1 ;
      RECT 5.21 0.33 5.4 2.63 ;
      RECT 4.315 2.44 5.4 2.63 ;
      RECT 8.24 1.9 9.135 2.09 ;
      RECT 3.925 1.99 4.22 2.18 ;
      RECT 5.68 2.085 7.515 2.275 ;
      RECT 0.2 0.33 0.39 2.77 ;
      RECT 0.2 2.58 4.115 2.77 ;
      RECT 3.925 1.99 4.115 3.02 ;
      RECT 7.325 2.085 7.515 3.04 ;
      RECT 5.68 1.275 5.87 3.02 ;
      RECT 3.925 2.83 5.87 3.02 ;
      RECT 8.24 1.9 8.43 3.04 ;
      RECT 7.325 2.85 8.43 3.04 ;
      RECT 7.81 0.325 8 1.7 ;
      RECT 6.49 1.5 8 1.69 ;
      RECT 7.76 1.51 10.04 1.7 ;
      RECT 7.76 1.5 7.95 2.62 ;
      RECT 7.715 2.425 7.995 2.62 ;
      RECT 9.425 0.35 9.615 0.795 ;
      RECT 11.045 0.51 11.235 0.795 ;
      RECT 9.425 0.605 11.235 0.795 ;
      RECT 8.525 0.51 8.715 1.31 ;
      RECT 8.525 1.12 10.43 1.31 ;
      RECT 10.24 1.12 10.43 2.205 ;
      RECT 11.69 1.715 11.88 2.205 ;
      RECT 9.555 2.015 11.88 2.205 ;
      RECT 9.555 2.015 9.84 2.54 ;
  END
END CLKLANAQV3_7TV50

MACRO CLKLANQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLANQV1_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.415 1.56 1.84 1.9 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.855 1.52 4.305 1.84 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.31 0.69 11.5 2.475 ;
        RECT 11.64 0.56 11.92 0.88 ;
        RECT 11.31 0.69 11.92 0.88 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.095 1.65 3.285 2.28 ;
        RECT 2.96 2 3.285 2.28 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 2.91 1.395 3.48 ;
        RECT 2.615 2.91 2.895 3.48 ;
        RECT 7.095 2.91 7.375 3.48 ;
        RECT 8.595 2.91 8.875 3.48 ;
        RECT 10.415 2.275 10.695 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.72 ;
        RECT 2.545 -0.12 2.825 0.72 ;
        RECT 4.405 -0.12 4.685 0.39 ;
        RECT 7.595 -0.12 7.875 0.735 ;
        RECT 10.785 -0.12 11.07 0.86 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 0.655 1.46 ;
        RECT -0.12 -0.24 12.6 1.32 ;
        RECT 8.7 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 0.655 1.32 8.7 3.94 ;
        RECT -0.58 1.46 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.49 0.455 3.68 0.78 ;
      RECT 5.04 0.455 5.23 0.78 ;
      RECT 3.49 0.59 5.23 0.78 ;
      RECT 2 0.455 2.19 1.17 ;
      RECT 0.68 0.98 5.65 1.17 ;
      RECT 2.115 0.98 2.305 2.29 ;
      RECT 2.025 2.1 2.305 2.29 ;
      RECT 5.94 0.935 8.25 1.125 ;
      RECT 5.94 0.455 6.13 2.32 ;
      RECT 5.045 2.13 6.13 2.32 ;
      RECT 6.33 1.325 6.61 1.515 ;
      RECT 0.2 0.455 0.39 2.71 ;
      RECT 4.595 1.65 4.785 2.71 ;
      RECT 6.33 1.325 6.53 2.71 ;
      RECT 0.2 2.52 9.265 2.71 ;
      RECT 9.075 2.52 9.265 2.93 ;
      RECT 8.54 0.455 8.73 1.57 ;
      RECT 7.07 1.325 8.73 1.515 ;
      RECT 8.095 1.38 10.16 1.57 ;
      RECT 8.095 1.325 8.285 2.32 ;
      RECT 8.005 2.13 8.285 2.32 ;
      RECT 9.085 0.625 10.575 0.815 ;
      RECT 10.385 0.625 10.575 1.995 ;
      RECT 9.55 1.805 11.07 1.995 ;
      RECT 9.55 1.805 9.74 2.475 ;
  END
END CLKLANQV1_7TV50

MACRO CLKLANQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLANQV2_7TV50 0 0 ;
  SIZE 12.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.415 1.56 1.84 1.9 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.855 1.52 4.305 1.84 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.31 0.56 11.5 2.895 ;
        RECT 11.31 0.56 11.92 0.88 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.095 1.65 3.285 2.28 ;
        RECT 2.96 2 3.285 2.28 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 2.91 1.395 3.48 ;
        RECT 2.615 2.91 2.895 3.48 ;
        RECT 7.095 2.91 7.375 3.48 ;
        RECT 8.595 2.91 8.875 3.48 ;
        RECT 10.415 2.275 10.695 3.48 ;
        RECT 8.595 3.235 10.695 3.48 ;
        RECT 12.115 2.32 12.395 3.48 ;
        RECT 0 3.24 12.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.72 ;
        RECT 1.055 -0.12 2.825 0.125 ;
        RECT 2.545 -0.12 2.825 0.72 ;
        RECT 4.405 -0.12 4.685 0.39 ;
        RECT 7.595 -0.12 7.875 0.735 ;
        RECT 10.785 -0.12 11.07 0.86 ;
        RECT 0 -0.12 12.96 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 0.655 1.46 ;
        RECT -0.12 -0.24 13.08 1.32 ;
        RECT 8.7 -0.24 13.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 0.655 1.32 8.7 3.94 ;
        RECT -0.58 1.46 13.54 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.49 0.455 3.68 0.78 ;
      RECT 5.04 0.455 5.23 0.78 ;
      RECT 3.49 0.59 5.23 0.78 ;
      RECT 2 0.455 2.19 1.17 ;
      RECT 0.68 0.98 5.65 1.17 ;
      RECT 2.115 0.98 2.305 2.29 ;
      RECT 2.025 2.1 2.305 2.29 ;
      RECT 5.94 0.935 8.25 1.125 ;
      RECT 5.94 0.455 6.13 2.32 ;
      RECT 5.045 2.13 6.13 2.32 ;
      RECT 6.42 1.325 6.7 1.515 ;
      RECT 0.2 0.435 0.39 2.71 ;
      RECT 4.595 1.65 4.785 2.71 ;
      RECT 6.42 1.325 6.62 2.71 ;
      RECT 9.075 1.76 9.265 2.71 ;
      RECT 0.2 2.52 9.265 2.71 ;
      RECT 8.54 0.455 8.73 1.515 ;
      RECT 7.22 1.325 10.16 1.515 ;
      RECT 9.88 1.325 10.16 1.685 ;
      RECT 8.095 1.325 8.285 2.32 ;
      RECT 8.005 2.13 8.285 2.32 ;
      RECT 9.085 0.5 10.575 0.69 ;
      RECT 10.385 1.805 11.07 1.995 ;
      RECT 10.385 0.5 10.575 2.075 ;
      RECT 9.55 1.885 10.575 2.075 ;
      RECT 9.55 1.885 9.74 2.475 ;
  END
END CLKLANQV2_7TV50

MACRO CLKLANQV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKLANQV3_7TV50 0 0 ;
  SIZE 13.44 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 1.415 1.56 1.84 1.9 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.855 1.52 4.305 1.84 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.31 1.465 11.5 2.475 ;
        RECT 11.6 0.58 11.92 0.845 ;
        RECT 11.73 0.58 11.92 1.655 ;
        RECT 11.31 1.465 13.2 1.655 ;
        RECT 13.01 1.465 13.2 2.475 ;
    END
  END Q
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.095 1.65 3.285 2.28 ;
        RECT 2.96 2 3.285 2.28 ;
    END
  END TE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 2.91 1.395 3.48 ;
        RECT 2.615 2.91 2.895 3.48 ;
        RECT 7.095 2.91 7.375 3.48 ;
        RECT 8.595 2.91 8.875 3.48 ;
        RECT 10.415 2.275 10.695 3.48 ;
        RECT 8.595 3.235 10.695 3.48 ;
        RECT 12.115 2.32 12.395 3.48 ;
        RECT 0 3.24 13.44 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.72 ;
        RECT 1.055 -0.12 2.825 0.125 ;
        RECT 2.545 -0.12 2.825 0.72 ;
        RECT 4.405 -0.12 4.685 0.39 ;
        RECT 7.595 -0.12 7.875 0.735 ;
        RECT 10.785 -0.12 11.07 0.86 ;
        RECT 12.585 -0.12 12.865 0.815 ;
        RECT 0 -0.12 13.44 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 0.655 1.46 ;
        RECT -0.12 -0.24 13.56 1.32 ;
        RECT 8.7 -0.24 13.56 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 0.655 1.32 8.7 3.94 ;
        RECT -0.58 1.46 14.02 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.49 0.455 3.68 0.78 ;
      RECT 5.04 0.455 5.23 0.78 ;
      RECT 3.49 0.59 5.23 0.78 ;
      RECT 2 0.455 2.19 1.17 ;
      RECT 0.68 0.98 5.65 1.17 ;
      RECT 2.115 0.98 2.305 2.29 ;
      RECT 2.025 2.1 2.305 2.29 ;
      RECT 5.94 0.935 8.25 1.125 ;
      RECT 5.94 0.455 6.13 2.32 ;
      RECT 5.045 2.13 6.13 2.32 ;
      RECT 6.42 1.325 6.7 1.515 ;
      RECT 0.2 0.435 0.39 2.71 ;
      RECT 4.595 1.65 4.785 2.71 ;
      RECT 6.42 1.325 6.62 2.71 ;
      RECT 9.075 1.76 9.265 2.71 ;
      RECT 0.2 2.52 9.265 2.71 ;
      RECT 8.54 0.455 8.73 1.515 ;
      RECT 7.07 1.325 10.16 1.515 ;
      RECT 9.88 1.325 10.16 1.685 ;
      RECT 8.095 1.325 8.285 2.32 ;
      RECT 8.005 2.13 8.285 2.32 ;
      RECT 9.085 0.5 10.575 0.69 ;
      RECT 10.385 1.805 11.07 1.995 ;
      RECT 10.385 0.5 10.575 2.075 ;
      RECT 9.55 1.885 10.575 2.075 ;
      RECT 9.55 1.885 9.74 2.475 ;
  END
END CLKLANQV3_7TV50

MACRO CLKMUX2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMUX2V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.87 1.425 4.445 1.8 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.345 1.52 1.815 1.85 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.08 1.36 1.32 ;
        RECT 0.83 1.125 2.51 1.32 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.545 1.485 3.48 ;
        RECT 4.455 2.545 4.735 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.815 ;
        RECT 4.455 -0.12 4.735 0.815 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 0.56 5.59 2.58 ;
        RECT 5.31 2.39 5.59 2.58 ;
        RECT 5.4 1.52 5.64 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.71 1.06 3.5 1.25 ;
      RECT 0.2 0.58 0.39 2.24 ;
      RECT 2.38 2 2.9 2.24 ;
      RECT 2.71 1.06 2.9 2.24 ;
      RECT 0.2 2.05 2.9 2.24 ;
      RECT 0.4 2.05 0.59 2.67 ;
      RECT 2.755 0.625 4.14 0.815 ;
      RECT 3.95 0.625 4.14 1.205 ;
      RECT 3.95 1.015 5.065 1.205 ;
      RECT 4.875 1.015 5.065 2.19 ;
      RECT 3.1 2 5.065 2.19 ;
      RECT 3.1 2 3.29 2.73 ;
      RECT 2.805 2.54 3.29 2.73 ;
  END
END CLKMUX2V1_7TV50

MACRO CLKMUX2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMUX2V2_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.455 1.47 1.875 1.815 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.855 1.56 4.42 1.815 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.75 2.025 0.94 2.415 ;
        RECT 3 1.075 3.245 2.415 ;
        RECT 0.75 2.225 3.245 2.415 ;
        RECT 3 1.075 3.435 1.27 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.095 2.775 1.375 3.48 ;
        RECT 4.43 2.795 4.71 3.48 ;
        RECT 6.255 2.405 6.535 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.08 -0.12 1.36 0.83 ;
        RECT 4.54 -0.12 4.82 0.58 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.52 5.735 1.84 ;
        RECT 5.545 0.595 5.735 2.52 ;
        RECT 5.405 2.33 5.735 2.52 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.225 1.08 2.67 1.27 ;
      RECT 0.225 0.595 0.415 2.695 ;
      RECT 0.225 2.505 0.505 2.695 ;
      RECT 2.78 0.64 4.255 0.83 ;
      RECT 4.065 0.64 4.255 1.27 ;
      RECT 4.065 1.08 5.255 1.27 ;
      RECT 4.62 1.08 4.81 2.595 ;
      RECT 3.865 2.405 4.81 2.595 ;
      RECT 3.865 2.405 4.055 2.94 ;
      RECT 2.83 2.75 4.055 2.94 ;
  END
END CLKMUX2V2_7TV50

MACRO CLKNAND2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKNAND2V1_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.56 1.865 1.98 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.12 1.52 0.36 1.86 ;
        RECT 0.12 1.67 0.87 1.86 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 2.4 0.495 3.48 ;
        RECT 1.915 2.4 2.195 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.12 0.445 0.74 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.11 0.64 1.3 2.475 ;
        RECT 1.08 1.04 1.32 1.36 ;
        RECT 1.11 0.64 2.145 0.83 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
END CLKNAND2V1_7TV50

MACRO CLKNAND2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKNAND2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.305 1.5 2.765 1.87 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.56 1.93 1.915 ;
        RECT 0.625 1.725 1.93 1.915 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.405 0.435 3.48 ;
        RECT 1.955 2.795 2.235 3.48 ;
        RECT 3.655 2.405 3.935 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.715 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.915 0.71 3.24 0.9 ;
        RECT 3 0.71 3.24 1.36 ;
        RECT 3.05 0.71 3.24 2.595 ;
        RECT 1.105 2.405 3.24 2.595 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.41 -0.24 3.705 1.53 ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.41 3.94 ;
        RECT 3.705 1.46 4.9 3.94 ;
        RECT -0.58 1.53 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2 0.32 4.11 0.51 ;
      RECT 3.92 0.32 4.11 0.76 ;
      RECT 0.2 0.57 0.39 1.105 ;
      RECT 2 0.32 2.195 1.105 ;
      RECT 0.2 0.915 2.195 1.105 ;
  END
END CLKNAND2V2_7TV50

MACRO CLKNAND2V3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKNAND2V3_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 1.52 3.72 2.11 ;
        RECT 3.265 1.83 3.72 2.11 ;
        RECT 4.015 1.83 4.205 2.11 ;
        RECT 3.265 1.92 4.205 2.11 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.52 2.28 2.065 ;
        RECT 1.435 1.875 2.65 2.065 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.405 0.475 3.48 ;
        RECT 1.895 2.795 2.175 3.48 ;
        RECT 3.595 2.795 3.875 3.48 ;
        RECT 5.295 2.405 5.575 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.845 -0.12 2.125 0.565 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.705 0.71 3.985 1.175 ;
        RECT 3.705 0.985 4.68 1.175 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.49 0.985 4.68 2.595 ;
        RECT 1.045 2.405 4.68 2.595 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.035 -0.24 4.475 1.53 ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.035 3.94 ;
        RECT 4.475 1.46 6.34 3.94 ;
        RECT -0.58 1.53 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.79 0.32 4.9 0.51 ;
      RECT 4.71 0.32 4.9 0.61 ;
      RECT 0.99 0.595 1.18 0.955 ;
      RECT 2.79 0.32 2.98 0.955 ;
      RECT 0.99 0.765 2.98 0.955 ;
  END
END CLKNAND2V3_7TV50

MACRO CLKNOR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKNOR2V1_7TV50 0 0 ;
  SIZE 2.88 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 2.045 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 0.88 1.8 ;
        RECT 0.82 1.61 1.01 2.04 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.4 2.355 0.68 3.48 ;
        RECT 0 3.24 2.88 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.29 -0.12 0.57 0.875 ;
        RECT 2.445 -0.12 2.725 0.83 ;
        RECT 0 -0.12 2.88 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.505 0.595 1.695 1.22 ;
        RECT 1.505 1.03 2.485 1.22 ;
        RECT 2 2.24 2.32 2.76 ;
        RECT 2.295 1.03 2.485 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.46 3.94 ;
    END
  END VNW
END CLKNOR2V1_7TV50

MACRO CLKNOR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKNOR2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 1.04 3.93 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.08 1.97 1.4 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.31 2.745 1.59 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.26 -0.12 1.54 0.815 ;
        RECT 3.06 -0.12 3.34 0.81 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.205 0.595 2.395 1.75 ;
        RECT 2.205 1.56 3.28 1.75 ;
        RECT 3.055 1.56 3.245 2.475 ;
        RECT 2.96 1.56 3.28 1.8 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.45 2.24 2.395 2.43 ;
      RECT 2.205 2.24 2.395 2.865 ;
      RECT 3.905 2.195 4.095 2.865 ;
      RECT 2.205 2.675 4.095 2.865 ;
  END
END CLKNOR2V2_7TV50

MACRO CLKNOR2V3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKNOR2V3_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.855 1.52 5.175 2.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.555 1.52 0.84 2.045 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.2 2.36 0.48 3.48 ;
        RECT 1.9 2.79 2.18 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.16 -0.12 2.44 0.59 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.305 0.6 1.495 1.195 ;
        RECT 1.305 1.005 3.79 1.195 ;
        RECT 3.385 1.52 3.79 1.84 ;
        RECT 3.6 0.6 3.79 2.435 ;
        RECT 3.6 2.245 5.595 2.435 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.98 -0.24 4.625 1.465 ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.98 3.94 ;
        RECT 4.625 1.46 6.34 3.94 ;
        RECT -0.58 1.465 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.05 2.345 2.985 2.54 ;
      RECT 2.795 2.345 2.985 2.925 ;
      RECT 2.795 2.735 4.73 2.925 ;
  END
END CLKNOR2V3_7TV50

MACRO CLKOR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKOR2V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.35 1.075 0.88 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.85 2.04 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.075 2.565 2.355 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.225 -0.12 0.505 0.875 ;
        RECT 2.025 -0.12 2.305 0.875 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.97 0.595 3.16 2.475 ;
        RECT 2.97 2 3.24 2.33 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.17 1.075 2.68 1.265 ;
      RECT 1.17 0.595 1.36 2.43 ;
      RECT 0.375 2.24 1.36 2.43 ;
  END
END CLKOR2V1_7TV50

MACRO CLKOR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKOR2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.42 1.52 0.9 1.86 ;
        RECT 0.615 1.52 0.9 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.465 1.495 1.745 1.995 ;
        RECT 1.395 1.495 1.84 1.84 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.94 2.745 2.22 3.48 ;
        RECT 3.79 2.3 4.07 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.19 -0.12 0.47 0.875 ;
        RECT 1.99 -0.12 2.27 0.83 ;
        RECT 1.99 -0.12 4.07 0.225 ;
        RECT 3.79 -0.12 4.07 0.78 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.935 0.595 3.125 2.475 ;
        RECT 2.935 1.07 3.28 1.385 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.135 0.595 1.325 1.265 ;
      RECT 1.135 1.075 2.67 1.265 ;
      RECT 2.04 1.075 2.23 2.43 ;
      RECT 0.24 2.24 2.23 2.43 ;
  END
END CLKOR2V2_7TV50

MACRO CLKOR2V3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKOR2V3_7TV50 0 0 ;
  SIZE 4.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.505 1.08 0.89 1.46 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.53 1.03 1.915 1.415 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.815 2.355 2.095 3.48 ;
        RECT 3.515 2.75 3.795 3.48 ;
        RECT 0 3.24 4.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 -0.12 0.475 0.875 ;
        RECT 1.995 -0.12 2.275 0.83 ;
        RECT 3.795 -0.12 4.075 0.875 ;
        RECT 0 -0.12 4.8 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.94 0.595 3.13 2.43 ;
        RECT 3.92 2.04 4.24 2.43 ;
        RECT 2.665 2.24 4.645 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.14 0.595 1.33 1.995 ;
      RECT 0.26 1.805 2.47 1.995 ;
      RECT 0.26 1.805 0.45 2.55 ;
  END
END CLKOR2V3_7TV50

MACRO CLKXOR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2V1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.08 3.28 1.32 ;
        RECT 2.77 1.13 5.075 1.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 1.52 4.355 2.04 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.555 2.925 0.835 3.48 ;
        RECT 4.405 2.655 4.685 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.4 0.875 ;
        RECT 4.405 -0.12 4.685 0.875 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.64 0.84 2.675 ;
        RECT 0.6 0.64 2.135 0.83 ;
        RECT 0.6 2.485 2.94 2.675 ;
        RECT 2.75 2.485 2.94 2.765 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.335 0.64 3.785 0.83 ;
      RECT 2.335 0.64 2.525 1.28 ;
      RECT 1.135 1.09 2.525 1.28 ;
      RECT 1.135 1.09 1.325 2.285 ;
      RECT 1.135 2.095 3.37 2.285 ;
      RECT 3.18 2.095 3.37 2.82 ;
      RECT 3.18 2.63 3.835 2.82 ;
      RECT 1.66 1.705 3.76 1.895 ;
      RECT 3.57 1.705 3.76 2.43 ;
      RECT 5.35 0.595 5.54 2.43 ;
      RECT 3.57 2.24 5.54 2.43 ;
  END
END CLKXOR2V1_7TV50

MACRO CLKXOR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2V2_7TV50 0 0 ;
  SIZE 8.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.445 1.745 7.725 2 ;
        RECT 7.48 1.56 8.08 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.535 1.52 1.065 1.8 ;
        RECT 0.77 1.52 1.065 2 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.385 2.36 0.665 3.48 ;
        RECT 2.21 2.795 2.49 3.48 ;
        RECT 6.11 2.245 6.39 3.48 ;
        RECT 7.82 2.405 8.1 3.48 ;
        RECT 0 3.24 8.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.44 0.76 ;
        RECT 2.195 -0.12 2.46 0.76 ;
        RECT 6.06 -0.12 6.345 0.715 ;
        RECT 8.1 -0.12 8.38 0.715 ;
        RECT 0 -0.12 8.64 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.055 0.725 4.335 1.35 ;
        RECT 4.055 1.08 4.8 1.35 ;
        RECT 4.61 1.08 4.8 1.69 ;
        RECT 4.61 1.5 5.87 1.69 ;
        RECT 5.68 1.5 5.87 2.55 ;
        RECT 4.76 2.36 5.87 2.55 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.805 -0.24 5.65 1.545 ;
        RECT -0.12 -0.24 8.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.805 3.94 ;
        RECT 5.65 1.46 9.22 3.94 ;
        RECT -0.58 1.545 9.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.155 0.725 3.435 0.915 ;
      RECT 3.245 0.725 3.435 2.55 ;
      RECT 3.155 2.36 3.435 2.55 ;
      RECT 3.635 1.115 3.825 2.08 ;
      RECT 3.635 1.89 5.43 2.08 ;
      RECT 2.765 0.32 5.19 0.51 ;
      RECT 5 0.32 5.19 0.96 ;
      RECT 1.23 0.48 1.42 1.17 ;
      RECT 1.23 0.98 2.955 1.17 ;
      RECT 1.335 2.395 2.955 2.585 ;
      RECT 2.765 0.32 2.955 2.985 ;
      RECT 2.765 2.795 5.9 2.985 ;
      RECT 5.495 0.545 5.685 1.14 ;
      RECT 7.125 0.48 7.315 1.14 ;
      RECT 5.495 0.95 7.315 1.14 ;
      RECT 7.015 0.95 7.205 2.48 ;
  END
END CLKXOR2V2_7TV50

MACRO CLKXOR2V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2V4_7TV50 0 0 ;
  SIZE 16.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.295 1.395 9.575 1.825 ;
        RECT 7.58 1.635 9.575 1.825 ;
        RECT 13.79 1.51 14.76 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4 1.56 3.46 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.405 0.435 3.48 ;
        RECT 1.855 2.405 2.135 3.48 ;
        RECT 3.555 2.405 3.835 3.48 ;
        RECT 12.485 2.795 12.765 3.48 ;
        RECT 14.185 2.795 14.465 3.48 ;
        RECT 15.885 2.405 16.165 3.48 ;
        RECT 0 3.24 16.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.755 -0.12 2.035 0.78 ;
        RECT 3.555 -0.12 3.835 0.83 ;
        RECT 12.38 -0.12 12.57 0.825 ;
        RECT 14.135 -0.12 14.415 0.78 ;
        RECT 0 -0.12 16.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.355 0.32 5.635 0.76 ;
        RECT 7.275 0.32 7.555 0.755 ;
        RECT 9.785 0.32 10.065 0.665 ;
        RECT 5.355 0.32 11.82 0.51 ;
        RECT 11.615 0.32 11.805 2.985 ;
        RECT 5.77 2.795 11.805 2.985 ;
        RECT 11.615 0.32 11.82 1.36 ;
        RECT 11.615 1.04 11.88 1.36 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 5.625 -0.24 12.185 1.535 ;
        RECT -0.12 -0.24 16.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.625 3.94 ;
        RECT 12.185 1.46 16.9 3.94 ;
        RECT -0.58 1.535 16.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.7 0.595 2.89 1.22 ;
      RECT 0.9 1.02 2.89 1.22 ;
      RECT 0.9 1.03 4.18 1.22 ;
      RECT 3.99 1.03 4.18 1.31 ;
      RECT 0.9 0.595 1.09 2.19 ;
      RECT 0.9 2 2.985 2.19 ;
      RECT 1.005 2 1.285 2.445 ;
      RECT 2.705 2 2.985 2.445 ;
      RECT 4.5 0.595 4.69 1.195 ;
      RECT 6.315 0.71 6.6 1.195 ;
      RECT 8.235 0.71 8.52 1.195 ;
      RECT 4.38 1.005 8.52 1.195 ;
      RECT 4.38 1.005 4.57 2.595 ;
      RECT 4.38 2.405 6.9 2.595 ;
      RECT 8.885 0.71 9.165 1.13 ;
      RECT 10.685 0.71 10.965 1.13 ;
      RECT 8.885 0.94 11 1.13 ;
      RECT 4.77 1.575 4.96 2.05 ;
      RECT 4.77 1.86 7.315 2.05 ;
      RECT 7.125 1.86 7.315 2.595 ;
      RECT 10.81 0.94 11 2.595 ;
      RECT 7.125 2.405 11 2.595 ;
      RECT 15.08 0.595 15.27 1.17 ;
      RECT 13.28 0.98 15.27 1.17 ;
      RECT 12.005 1.92 12.195 2.435 ;
      RECT 13.28 0.595 13.47 2.435 ;
      RECT 12.005 2.245 15.315 2.435 ;
  END
END CLKXOR2V4_7TV50

MACRO DEL1V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DEL1V1_7TV50 0 0 ;
  SIZE 4.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.94 1.47 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.675 1.345 3.48 ;
        RECT 3.515 2.55 3.795 3.48 ;
        RECT 0 3.24 4.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.83 ;
        RECT 3.465 -0.12 3.745 0.83 ;
        RECT 0 -0.12 4.8 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.41 0.595 4.6 2.475 ;
        RECT 4.41 1.52 4.68 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.805 1.71 1.995 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 2.01 0.595 2.2 2.475 ;
      RECT 2.01 1.44 2.92 1.63 ;
      RECT 2.01 1.44 2.21 2.475 ;
      RECT 2.6 0.595 2.79 1.22 ;
      RECT 2.6 1.03 3.595 1.22 ;
      RECT 3.405 1.03 3.595 2.305 ;
      RECT 2.66 2.115 3.595 2.305 ;
      RECT 2.66 2.115 2.85 2.475 ;
  END
END DEL1V1_7TV50

MACRO DEL1V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DEL1V2_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 1.04 1.09 1.43 ;
        RECT 0.72 1.04 1.32 1.36 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.18 2.25 1.46 3.48 ;
        RECT 3.58 2.25 3.86 3.48 ;
        RECT 5.285 2.795 5.565 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.13 -0.12 1.41 0.83 ;
        RECT 3.58 -0.12 3.86 0.83 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.48 0.595 4.67 2.43 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.435 0.595 4.715 0.91 ;
        RECT 4.435 2.16 4.715 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.215 0.595 0.405 1.995 ;
      RECT 0.215 1.805 1.845 1.995 ;
      RECT 0.315 1.805 0.505 2.475 ;
      RECT 2.135 1.48 2.575 1.67 ;
      RECT 2.135 0.595 2.325 2.475 ;
      RECT 2.725 0.595 2.915 1.28 ;
      RECT 2.775 1.805 4.235 1.995 ;
      RECT 2.775 1.09 2.965 2.475 ;
  END
END DEL1V2_7TV50

MACRO DEL2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DEL2V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.04 1.32 1.41 ;
        RECT 0.675 1.13 1.32 1.41 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.215 2.675 1.495 3.48 ;
        RECT 5.265 2.24 5.545 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.215 -0.12 1.495 0.83 ;
        RECT 5.325 -0.12 5.605 0.83 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.33 0.595 6.52 2.475 ;
        RECT 6.33 1.52 6.6 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.24 0.595 0.43 1.995 ;
      RECT 0.24 1.805 1.93 1.995 ;
      RECT 0.285 1.805 0.475 2.475 ;
      RECT 3.02 1.43 3.335 1.62 ;
      RECT 3.02 0.595 3.21 2.475 ;
      RECT 3.61 1.075 6.04 1.265 ;
      RECT 3.61 0.595 3.8 2.475 ;
  END
END DEL2V1_7TV50

MACRO DEL2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DEL2V2_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.875 1.56 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 2.3 1.355 3.48 ;
        RECT 5.065 2.3 5.345 3.48 ;
        RECT 6.765 2.795 7.045 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 -0.12 1.345 0.83 ;
        RECT 5.065 -0.12 5.345 0.83 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.96 1.52 6.15 2.475 ;
        RECT 6.01 0.595 6.2 1.71 ;
        RECT 5.96 1.52 6.6 1.71 ;
        RECT 6.36 1.52 6.6 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.21 1.805 1.79 1.995 ;
      RECT 0.21 0.595 0.4 2.475 ;
      RECT 2.82 1.485 3.135 1.675 ;
      RECT 2.82 0.595 3.01 2.475 ;
      RECT 3.41 1.485 5.24 1.675 ;
      RECT 3.41 0.595 3.6 2.475 ;
  END
END DEL2V2_7TV50

MACRO DEL4V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DEL4V1_7TV50 0 0 ;
  SIZE 9.6 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.04 1.8 1.365 ;
        RECT 0.865 1.175 1.8 1.365 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.1 2.32 1.38 3.48 ;
        RECT 8.165 2.265 8.445 3.48 ;
        RECT 0 3.24 9.6 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 -0.12 1.355 0.83 ;
        RECT 8.265 -0.12 8.545 0.83 ;
        RECT 0 -0.12 9.6 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.21 0.595 9.4 2.475 ;
        RECT 9.21 1.52 9.48 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.72 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 10.18 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.22 1.805 4.13 1.995 ;
      RECT 0.22 0.595 0.41 2.475 ;
      RECT 4.42 1.445 4.925 1.635 ;
      RECT 4.42 0.595 4.61 2.475 ;
      RECT 4.955 0.64 5.315 0.83 ;
      RECT 5.125 1.48 8.72 1.67 ;
      RECT 5.125 0.64 5.315 2.43 ;
      RECT 5 2.235 5.315 2.43 ;
  END
END DEL4V1_7TV50

MACRO DEL4V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DEL4V2_7TV50 0 0 ;
  SIZE 10.56 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.9 1.56 1.36 1.875 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.135 2.7 1.415 3.48 ;
        RECT 8.325 2.26 8.605 3.48 ;
        RECT 10.125 2.36 10.405 3.48 ;
        RECT 0 3.24 10.56 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.135 -0.12 1.415 0.875 ;
        RECT 8.325 -0.12 8.605 0.76 ;
        RECT 10.125 -0.12 10.405 0.805 ;
        RECT 0 -0.12 10.56 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.27 0.525 9.46 2.64 ;
        RECT 9.24 1.52 9.48 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 10.68 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 11.14 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.575 1.805 2.59 1.995 ;
      RECT 0.27 0.595 0.46 2.475 ;
      RECT 1.575 1.805 1.765 2.475 ;
      RECT 0.27 2.275 1.765 2.475 ;
      RECT 4.48 1.485 5.15 1.675 ;
      RECT 4.48 0.595 4.67 2.475 ;
      RECT 5.025 0.57 5.6 0.76 ;
      RECT 5.41 0.57 5.6 2.43 ;
      RECT 5.41 1.005 8.98 1.195 ;
      RECT 5.41 1.005 5.61 2.43 ;
      RECT 5.025 2.24 5.61 2.43 ;
  END
END DEL4V2_7TV50

MACRO DQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DQV1_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 1.12 1.36 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.95 1.56 3.425 1.87 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.065 0.595 12.255 2.475 ;
        RECT 12.065 1.52 12.36 1.84 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.135 2.925 1.365 3.48 ;
        RECT 2.67 2.305 2.95 3.48 ;
        RECT 5.985 2.925 6.265 3.48 ;
        RECT 9.63 2.39 9.91 3.48 ;
        RECT 11.17 2.285 11.45 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.07 -0.12 1.35 0.84 ;
        RECT 2.56 -0.12 2.84 0.935 ;
        RECT 6.07 -0.12 6.35 0.935 ;
        RECT 9.63 -0.12 9.91 0.77 ;
        RECT 11.12 -0.12 11.4 0.61 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.175 -0.24 8.575 1.57 ;
        RECT -0.12 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.175 3.94 ;
        RECT 8.575 1.46 13.06 3.94 ;
        RECT -0.58 1.57 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.17 0.64 0.45 0.83 ;
      RECT 0.17 1.815 1.835 2.005 ;
      RECT 0.17 0.64 0.36 2.54 ;
      RECT 0.17 2.35 0.46 2.54 ;
      RECT 1.97 0.64 2.265 0.83 ;
      RECT 2.075 1.17 4.125 1.36 ;
      RECT 3.845 1.17 4.125 1.41 ;
      RECT 2.075 0.64 2.265 2.585 ;
      RECT 4.36 0.42 4.55 1.375 ;
      RECT 4.36 1.185 6.725 1.375 ;
      RECT 4.37 1.185 4.56 2.585 ;
      RECT 5.55 1.915 7.205 2.105 ;
      RECT 7.015 0.705 7.205 2.585 ;
      RECT 4.845 1.87 5.035 2.645 ;
      RECT 4.845 2.455 6.735 2.645 ;
      RECT 6.545 2.455 6.735 3.01 ;
      RECT 7.445 1.85 7.635 3.01 ;
      RECT 6.545 2.82 7.635 3.01 ;
      RECT 7.495 1.185 8.445 1.375 ;
      RECT 8.255 1.185 8.445 2.36 ;
      RECT 7.87 0.745 8.935 0.935 ;
      RECT 8.745 1.625 10.135 1.815 ;
      RECT 8.745 0.745 8.935 2.75 ;
      RECT 7.835 2.56 8.935 2.75 ;
      RECT 9.19 1.075 11.775 1.265 ;
      RECT 10.575 0.565 10.765 2.48 ;
  END
END DQV1_7TV50

MACRO DQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DQV2_7TV50 0 0 ;
  SIZE 13.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.755 1.04 1.32 1.36 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.37 1.56 2.875 1.9 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.12 1.52 12.46 1.84 ;
        RECT 12.27 0.595 12.46 2.475 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.02 2.53 1.3 3.48 ;
        RECT 2.46 2.52 2.74 3.48 ;
        RECT 6.095 2.52 6.375 3.48 ;
        RECT 9.835 2.795 10.115 3.48 ;
        RECT 11.375 2.39 11.655 3.48 ;
        RECT 13.075 2.39 13.355 3.48 ;
        RECT 0 3.24 13.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.13 -0.12 1.41 0.83 ;
        RECT 2.62 -0.12 2.9 0.94 ;
        RECT 6.13 -0.12 6.41 0.94 ;
        RECT 9.835 -0.12 10.115 0.78 ;
        RECT 11.325 -0.12 11.605 0.635 ;
        RECT 13.125 -0.12 13.405 0.635 ;
        RECT 0 -0.12 13.92 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.175 -0.24 8.575 1.57 ;
        RECT -0.12 -0.24 14.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.175 3.94 ;
        RECT 8.575 1.46 14.5 3.94 ;
        RECT -0.58 1.57 14.5 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.23 0.64 0.515 0.83 ;
      RECT 0.23 0.64 0.42 2.72 ;
      RECT 0.23 2.095 1.675 2.285 ;
      RECT 0.23 2.095 0.425 2.72 ;
      RECT 0.17 2.53 0.45 2.72 ;
      RECT 2.075 0.595 2.265 1.36 ;
      RECT 1.915 1.17 3.395 1.36 ;
      RECT 3.205 1.17 3.395 2.105 ;
      RECT 3.205 1.915 3.82 2.105 ;
      RECT 3.63 1.87 3.82 2.15 ;
      RECT 1.915 1.17 2.105 2.765 ;
      RECT 4.42 1.185 6.835 1.375 ;
      RECT 4.42 0.675 4.61 2.585 ;
      RECT 7.075 0.705 7.265 1.93 ;
      RECT 5.71 1.74 7.265 1.93 ;
      RECT 7 1.74 7.19 2.585 ;
      RECT 3.975 1.14 4.21 1.42 ;
      RECT 5.015 2.13 6.765 2.32 ;
      RECT 4.02 1.14 4.21 2.975 ;
      RECT 6.575 2.13 6.765 3.01 ;
      RECT 5.015 1.87 5.205 2.975 ;
      RECT 4.02 2.785 5.205 2.975 ;
      RECT 7.505 1.85 7.695 3.01 ;
      RECT 6.575 2.82 7.695 3.01 ;
      RECT 7.555 1.185 8.61 1.375 ;
      RECT 8.42 1.185 8.61 2.36 ;
      RECT 7.93 0.75 9 0.94 ;
      RECT 8.81 1.81 10.49 2 ;
      RECT 8.81 0.75 9 2.75 ;
      RECT 7.915 2.56 9 2.75 ;
      RECT 10.78 0.565 10.97 1.265 ;
      RECT 9.42 1.075 11.98 1.265 ;
      RECT 10.73 1.075 10.92 2.48 ;
  END
END DQV2_7TV50

MACRO DRNQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DRNQV1_7TV50 0 0 ;
  SIZE 14.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.34 1.52 0.84 1.84 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.535 3.055 1.815 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.01 0.58 14.2 2.435 ;
        RECT 13.675 2.245 14.2 2.435 ;
        RECT 14.01 1.52 14.28 1.84 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.36 1.56 6 1.8 ;
        RECT 5.81 1.56 6 2.155 ;
        RECT 5.81 1.965 7.07 2.155 ;
        RECT 6.88 1.965 7.07 2.53 ;
        RECT 6.88 2.34 8.04 2.53 ;
        RECT 7.85 2.34 8.04 2.97 ;
        RECT 10.735 1.725 10.925 2.97 ;
        RECT 7.85 2.78 10.925 2.97 ;
        RECT 10.735 1.725 11.78 1.915 ;
    END
  END RDN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.355 0.435 3.48 ;
        RECT 2.445 2.355 2.725 3.48 ;
        RECT 5.81 2.745 6.09 3.48 ;
        RECT 7.37 2.73 7.65 3.48 ;
        RECT 11.125 2.405 11.405 3.48 ;
        RECT 12.825 2.405 13.105 3.48 ;
        RECT 0 3.24 14.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.835 ;
        RECT 2.57 -0.12 2.85 0.945 ;
        RECT 7.035 -0.12 7.315 0.715 ;
        RECT 10.775 -0.12 11.055 0.7 ;
        RECT 13.065 -0.12 13.345 0.565 ;
        RECT 0 -0.12 14.4 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.38 -0.24 10.41 1.575 ;
        RECT -0.12 -0.24 14.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.12 3.94 ;
        RECT 10.41 1.46 14.98 3.94 ;
        RECT -0.58 1.575 14.98 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.055 0.64 1.44 0.83 ;
      RECT 1.25 0.64 1.44 2.545 ;
      RECT 1.005 2.355 1.44 2.545 ;
      RECT 1.69 1.145 3.905 1.335 ;
      RECT 3.715 1.145 3.905 2.16 ;
      RECT 1.69 0.71 1.88 2.59 ;
      RECT 1.64 2.31 1.88 2.59 ;
      RECT 4.895 2.355 6.68 2.545 ;
      RECT 4.315 1.17 7.93 1.36 ;
      RECT 7.65 1.17 7.93 1.38 ;
      RECT 4.315 0.71 4.505 2.545 ;
      RECT 4.045 2.355 4.505 2.545 ;
      RECT 6.935 1.56 7.41 1.75 ;
      RECT 8.16 0.71 8.35 1.805 ;
      RECT 7.22 1.615 8.445 1.805 ;
      RECT 8.255 1.615 8.445 2.545 ;
      RECT 8.255 2.355 8.56 2.545 ;
      RECT 8.685 1.145 8.875 2.11 ;
      RECT 8.685 1.92 10.105 2.11 ;
      RECT 9.015 0.755 10.12 0.945 ;
      RECT 9.93 0.755 10.12 1.535 ;
      RECT 9.93 1.335 12.45 1.525 ;
      RECT 9.93 1.335 10.515 1.535 ;
      RECT 10.315 1.335 10.515 2.545 ;
      RECT 9.305 2.355 10.515 2.545 ;
      RECT 12.52 0.465 12.71 1.135 ;
      RECT 10.4 0.94 12.71 1.135 ;
      RECT 10.4 0.945 13.535 1.135 ;
      RECT 13.345 0.945 13.535 2.035 ;
      RECT 12.02 1.845 13.535 2.035 ;
      RECT 12.02 1.845 12.21 2.48 ;
  END
END DRNQV1_7TV50

MACRO DRNQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DRNQV2_7TV50 0 0 ;
  SIZE 15.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.34 1.52 0.84 1.84 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.535 3.055 1.815 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.01 0.525 14.2 2.435 ;
        RECT 13.675 2.245 14.2 2.435 ;
        RECT 14.01 1.52 14.28 1.84 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.36 1.56 6 1.8 ;
        RECT 5.81 1.56 6 2.155 ;
        RECT 5.81 1.965 7.07 2.155 ;
        RECT 6.88 1.965 7.07 2.53 ;
        RECT 6.88 2.34 8.04 2.53 ;
        RECT 7.85 2.34 8.04 2.97 ;
        RECT 10.735 1.725 10.925 2.97 ;
        RECT 7.85 2.78 10.925 2.97 ;
        RECT 10.735 1.725 11.78 1.915 ;
    END
  END RDN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.355 0.435 3.48 ;
        RECT 2.445 2.355 2.725 3.48 ;
        RECT 5.81 2.745 6.09 3.48 ;
        RECT 7.37 2.73 7.65 3.48 ;
        RECT 11.125 2.405 11.405 3.48 ;
        RECT 12.825 2.405 13.105 3.48 ;
        RECT 14.525 2.405 14.805 3.48 ;
        RECT 0 3.24 15.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.835 ;
        RECT 2.57 -0.12 2.85 0.945 ;
        RECT 7.035 -0.12 7.315 0.715 ;
        RECT 10.775 -0.12 11.055 0.7 ;
        RECT 13.065 -0.12 13.345 0.565 ;
        RECT 14.865 -0.12 15.145 0.57 ;
        RECT 0 -0.12 15.36 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.38 -0.24 10.41 1.575 ;
        RECT -0.12 -0.24 15.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.12 3.94 ;
        RECT 10.41 1.46 15.94 3.94 ;
        RECT -0.58 1.575 15.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.055 0.64 1.44 0.83 ;
      RECT 1.25 0.64 1.44 2.545 ;
      RECT 1.005 2.355 1.44 2.545 ;
      RECT 1.69 1.145 3.905 1.335 ;
      RECT 3.715 1.145 3.905 2.16 ;
      RECT 1.69 0.71 1.88 2.59 ;
      RECT 1.64 2.31 1.88 2.59 ;
      RECT 4.895 2.355 6.68 2.545 ;
      RECT 4.315 1.17 7.93 1.36 ;
      RECT 7.65 1.17 7.93 1.38 ;
      RECT 4.315 0.71 4.505 2.545 ;
      RECT 4.045 2.355 4.505 2.545 ;
      RECT 6.935 1.56 7.41 1.75 ;
      RECT 8.16 0.71 8.35 1.805 ;
      RECT 7.22 1.615 8.445 1.805 ;
      RECT 8.255 1.615 8.445 2.545 ;
      RECT 8.255 2.355 8.56 2.545 ;
      RECT 8.685 1.145 8.875 2.11 ;
      RECT 8.685 1.92 10.105 2.11 ;
      RECT 9.015 0.755 10.12 0.945 ;
      RECT 9.93 0.755 10.12 1.535 ;
      RECT 9.93 1.335 12.45 1.525 ;
      RECT 9.93 1.335 10.515 1.535 ;
      RECT 10.315 1.335 10.515 2.545 ;
      RECT 9.305 2.355 10.515 2.545 ;
      RECT 12.52 0.465 12.71 1.135 ;
      RECT 10.4 0.94 12.71 1.135 ;
      RECT 10.4 0.945 13.535 1.135 ;
      RECT 13.345 0.945 13.535 2.035 ;
      RECT 12.02 1.845 13.535 2.035 ;
      RECT 12.02 1.845 12.21 2.48 ;
  END
END DRNQV2_7TV50

MACRO DRQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DRQV1_7TV50 0 0 ;
  SIZE 14.88 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.8 1.04 1.36 1.32 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.37 1.56 2.875 1.85 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.465 0.595 14.655 2.475 ;
        RECT 14.465 1.52 14.76 1.845 ;
    END
  END Q
  PIN RD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.11 1.075 11.44 1.32 ;
        RECT 11.11 1.075 11.785 1.265 ;
    END
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.02 2.35 1.3 3.48 ;
        RECT 2.46 2.305 2.74 3.48 ;
        RECT 6.035 2.925 6.27 3.48 ;
        RECT 11.84 2.305 12.12 3.48 ;
        RECT 13.57 2.39 13.85 3.48 ;
        RECT 0 3.24 14.88 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.13 -0.12 1.41 0.84 ;
        RECT 2.62 -0.12 2.9 0.94 ;
        RECT 6.02 -0.12 6.3 0.94 ;
        RECT 7.88 -0.12 8.16 0.615 ;
        RECT 11.13 -0.12 11.41 0.83 ;
        RECT 13.52 -0.12 13.805 0.83 ;
        RECT 0 -0.12 14.88 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.255 -0.24 10.015 1.57 ;
        RECT -0.12 -0.24 15 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.255 3.94 ;
        RECT 10.015 1.46 15.46 3.94 ;
        RECT -0.58 1.57 15.46 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.23 0.64 0.515 0.83 ;
      RECT 0.23 0.64 0.43 2.105 ;
      RECT 0.23 1.915 1.675 2.105 ;
      RECT 0.23 0.64 0.425 2.54 ;
      RECT 0.17 2.35 0.45 2.54 ;
      RECT 2.075 0.595 2.265 1.36 ;
      RECT 1.915 1.17 3.395 1.36 ;
      RECT 3.205 1.17 3.395 2.06 ;
      RECT 3.205 1.87 3.82 2.06 ;
      RECT 3.63 1.87 3.82 2.15 ;
      RECT 1.915 1.17 2.105 2.585 ;
      RECT 4.32 0.75 4.61 0.94 ;
      RECT 4.42 1.445 7.455 1.635 ;
      RECT 7.265 1.445 7.455 2.15 ;
      RECT 4.42 0.75 4.61 2.585 ;
      RECT 6.92 0.75 7.34 0.94 ;
      RECT 8.33 0.75 8.75 0.94 ;
      RECT 7.15 0.815 8.52 1.005 ;
      RECT 5.6 1.915 7.05 2.105 ;
      RECT 6.86 1.915 7.05 2.54 ;
      RECT 7.655 0.815 7.845 2.54 ;
      RECT 6.86 2.35 8.92 2.54 ;
      RECT 3.92 1.14 4.21 1.42 ;
      RECT 4.895 2.535 6.66 2.725 ;
      RECT 6.47 2.535 6.66 2.93 ;
      RECT 4.02 1.14 4.21 2.975 ;
      RECT 9.145 1.87 9.335 2.93 ;
      RECT 6.47 2.74 9.335 2.93 ;
      RECT 4.895 1.87 5.085 2.975 ;
      RECT 4.02 2.785 5.085 2.975 ;
      RECT 8.925 1.185 10.1 1.375 ;
      RECT 9.91 1.185 10.1 2.15 ;
      RECT 9.37 0.75 10.49 0.94 ;
      RECT 12.075 0.595 12.265 1.71 ;
      RECT 10.3 1.52 13.375 1.71 ;
      RECT 10.3 0.75 10.49 2.54 ;
      RECT 9.535 2.35 10.49 2.54 ;
      RECT 9.535 2.305 9.725 2.585 ;
      RECT 12.665 0.595 12.855 1.22 ;
      RECT 12.665 1.03 14.13 1.22 ;
      RECT 13.94 1.03 14.13 2.1 ;
      RECT 10.715 1.91 14.13 2.1 ;
      RECT 12.765 1.91 12.955 2.475 ;
  END
END DRQV1_7TV50

MACRO DRQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DRQV2_7TV50 0 0 ;
  SIZE 15.84 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.8 1.04 1.36 1.32 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.37 1.56 2.875 1.85 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.465 0.595 14.655 2.475 ;
        RECT 14.465 1.52 14.76 1.845 ;
    END
  END Q
  PIN RD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.11 1.075 11.44 1.32 ;
        RECT 11.11 1.075 11.785 1.265 ;
    END
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.02 2.35 1.3 3.48 ;
        RECT 2.46 2.305 2.74 3.48 ;
        RECT 6.035 2.925 6.27 3.48 ;
        RECT 11.84 2.305 12.12 3.48 ;
        RECT 13.57 2.39 13.85 3.48 ;
        RECT 15.27 2.39 15.55 3.48 ;
        RECT 0 3.24 15.84 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.13 -0.12 1.41 0.84 ;
        RECT 2.62 -0.12 2.9 0.94 ;
        RECT 6.02 -0.12 6.3 0.94 ;
        RECT 7.88 -0.12 8.16 0.615 ;
        RECT 11.13 -0.12 11.41 0.83 ;
        RECT 13.52 -0.12 13.805 0.83 ;
        RECT 15.315 -0.12 15.6 0.83 ;
        RECT 0 -0.12 15.84 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.255 -0.24 10.015 1.57 ;
        RECT -0.12 -0.24 15.96 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.255 3.94 ;
        RECT 10.015 1.46 16.42 3.94 ;
        RECT -0.58 1.57 16.42 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.23 0.64 0.515 0.83 ;
      RECT 0.23 0.64 0.43 2.105 ;
      RECT 0.23 1.915 1.675 2.105 ;
      RECT 0.23 0.64 0.425 2.54 ;
      RECT 0.17 2.35 0.45 2.54 ;
      RECT 2.075 0.595 2.265 1.36 ;
      RECT 1.915 1.17 3.395 1.36 ;
      RECT 3.205 1.17 3.395 2.06 ;
      RECT 3.205 1.87 3.82 2.06 ;
      RECT 3.63 1.87 3.82 2.15 ;
      RECT 1.915 1.17 2.105 2.585 ;
      RECT 4.32 0.75 4.61 0.94 ;
      RECT 4.42 1.445 7.455 1.635 ;
      RECT 7.265 1.445 7.455 2.15 ;
      RECT 4.42 0.75 4.61 2.585 ;
      RECT 6.92 0.75 7.34 0.94 ;
      RECT 8.33 0.75 8.75 0.94 ;
      RECT 7.15 0.815 8.52 1.005 ;
      RECT 5.6 1.915 7.05 2.105 ;
      RECT 6.86 1.915 7.05 2.54 ;
      RECT 7.655 0.815 7.845 2.54 ;
      RECT 6.86 2.35 8.92 2.54 ;
      RECT 3.92 1.14 4.21 1.42 ;
      RECT 4.895 2.535 6.66 2.725 ;
      RECT 6.47 2.535 6.66 2.93 ;
      RECT 4.02 1.14 4.21 2.975 ;
      RECT 9.145 1.87 9.335 2.93 ;
      RECT 6.47 2.74 9.335 2.93 ;
      RECT 4.895 1.87 5.085 2.975 ;
      RECT 4.02 2.785 5.085 2.975 ;
      RECT 8.925 1.185 10.1 1.375 ;
      RECT 9.91 1.185 10.1 2.15 ;
      RECT 9.37 0.75 10.49 0.94 ;
      RECT 12.075 0.595 12.265 1.71 ;
      RECT 10.3 1.52 13.375 1.71 ;
      RECT 10.3 0.75 10.49 2.54 ;
      RECT 9.535 2.35 10.49 2.54 ;
      RECT 9.535 2.305 9.725 2.585 ;
      RECT 12.665 0.595 12.855 1.22 ;
      RECT 12.665 1.03 14.13 1.22 ;
      RECT 13.94 1.03 14.13 2.1 ;
      RECT 10.715 1.91 14.13 2.1 ;
      RECT 12.765 1.91 12.955 2.475 ;
  END
END DRQV2_7TV50

MACRO DSRNQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DSRNQV1_7TV50 0 0 ;
  SIZE 17.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.875 1 1.32 1.385 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.24 0.785 3.43 1.32 ;
        RECT 2.96 1.08 3.43 1.32 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.75 0.58 16.94 2.76 ;
        RECT 16.27 2.52 16.94 2.76 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.095 2.04 8.285 2.675 ;
        RECT 5.8 2.485 8.285 2.675 ;
        RECT 8.095 2.04 8.56 2.28 ;
        RECT 8.095 2.09 9.405 2.28 ;
        RECT 9.215 2.09 9.405 2.885 ;
        RECT 9.215 2.695 15.195 2.885 ;
    END
  END RDN
  PIN SDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.475 1.08 10.665 1.83 ;
        RECT 10.475 1.08 10.96 1.32 ;
        RECT 10.475 1.08 12.47 1.27 ;
    END
  END SDN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.38 2.24 1.66 3.48 ;
        RECT 2.82 2.26 3.1 3.48 ;
        RECT 8.615 2.615 8.895 3.48 ;
        RECT 15.45 2.615 15.73 3.48 ;
        RECT 0 3.24 17.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.33 -0.12 1.61 0.765 ;
        RECT 2.82 -0.12 3.1 0.57 ;
        RECT 7.79 -0.12 8.025 0.61 ;
        RECT 13.515 -0.12 13.795 0.625 ;
        RECT 15.805 -0.12 16.085 0.6 ;
        RECT 0 -0.12 17.28 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.935 1.46 ;
        RECT -0.12 -0.24 17.4 1.25 ;
        RECT 11.9 -0.24 17.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.935 1.25 11.9 3.94 ;
        RECT -0.58 1.46 17.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.475 0.52 0.665 1.99 ;
      RECT 0.475 1.8 2.035 1.99 ;
      RECT 0.575 1.8 0.765 2.475 ;
      RECT 5.33 2.03 7.325 2.22 ;
      RECT 4.465 0.375 7.59 0.565 ;
      RECT 7.4 0.375 7.59 1.05 ;
      RECT 7.4 0.86 8.475 1.05 ;
      RECT 4.465 0.375 4.655 2.485 ;
      RECT 4.94 0.83 7.2 1.02 ;
      RECT 7.01 0.83 7.2 1.44 ;
      RECT 9.695 0.89 9.885 1.44 ;
      RECT 7.01 1.25 9.885 1.44 ;
      RECT 2.275 1.815 4.225 2.005 ;
      RECT 2.275 0.53 2.465 2.49 ;
      RECT 3.755 1.815 3.945 2.875 ;
      RECT 4.94 0.83 5.13 2.875 ;
      RECT 3.755 2.685 5.13 2.875 ;
      RECT 9.41 0.425 10.395 0.62 ;
      RECT 6.615 1.55 6.805 1.83 ;
      RECT 10.085 0.425 10.275 1.83 ;
      RECT 6.615 1.64 10.275 1.83 ;
      RECT 9.63 1.64 9.82 2.265 ;
      RECT 7.68 1.64 7.87 2.285 ;
      RECT 11.46 2.26 13.16 2.45 ;
      RECT 11.015 0.43 12.95 0.62 ;
      RECT 12.76 0.955 14.385 1.145 ;
      RECT 12.76 0.43 12.95 1.99 ;
      RECT 10.91 1.8 12.95 1.99 ;
      RECT 10.91 1.8 11.1 2.45 ;
      RECT 10.555 2.26 11.1 2.45 ;
      RECT 14.1 0.43 14.775 0.62 ;
      RECT 13.35 1.79 16.125 1.98 ;
      RECT 14.585 0.43 14.775 2.475 ;
  END
END DSRNQV1_7TV50

MACRO DSRNQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DSRNQV2_7TV50 0 0 ;
  SIZE 18.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.875 1 1.32 1.385 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.24 0.785 3.43 1.32 ;
        RECT 2.96 1.08 3.43 1.32 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.75 0.58 16.94 2.76 ;
        RECT 16.27 2.52 16.94 2.76 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.095 2.04 8.285 2.675 ;
        RECT 5.8 2.485 8.285 2.675 ;
        RECT 8.095 2.04 8.56 2.28 ;
        RECT 8.095 2.09 9.405 2.28 ;
        RECT 9.215 2.09 9.405 2.885 ;
        RECT 9.215 2.695 15.195 2.885 ;
    END
  END RDN
  PIN SDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.475 1.08 10.665 1.83 ;
        RECT 10.475 1.08 10.96 1.32 ;
        RECT 10.475 1.08 12.47 1.27 ;
    END
  END SDN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.38 2.24 1.66 3.48 ;
        RECT 2.82 2.26 3.1 3.48 ;
        RECT 8.615 2.615 8.895 3.48 ;
        RECT 15.45 2.615 15.73 3.48 ;
        RECT 17.15 2.395 17.43 3.48 ;
        RECT 0 3.24 18.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.33 -0.12 1.61 0.765 ;
        RECT 2.82 -0.12 3.1 0.57 ;
        RECT 7.79 -0.12 8.025 0.61 ;
        RECT 13.515 -0.12 13.795 0.625 ;
        RECT 15.805 -0.12 16.085 0.6 ;
        RECT 17.605 -0.12 17.885 0.73 ;
        RECT 0 -0.12 18.24 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.935 1.46 ;
        RECT -0.12 -0.24 18.36 1.25 ;
        RECT 11.9 -0.24 18.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.935 1.25 11.9 3.94 ;
        RECT -0.58 1.46 18.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.475 0.52 0.665 1.99 ;
      RECT 0.475 1.8 2.035 1.99 ;
      RECT 0.575 1.8 0.765 2.475 ;
      RECT 5.33 2.03 7.325 2.22 ;
      RECT 4.465 0.375 7.59 0.565 ;
      RECT 7.4 0.375 7.59 1.05 ;
      RECT 7.4 0.86 8.475 1.05 ;
      RECT 4.465 0.375 4.655 2.485 ;
      RECT 4.94 0.83 7.2 1.02 ;
      RECT 7.01 0.83 7.2 1.44 ;
      RECT 9.695 0.89 9.885 1.44 ;
      RECT 7.01 1.25 9.885 1.44 ;
      RECT 2.275 1.815 4.225 2.005 ;
      RECT 2.275 0.53 2.465 2.49 ;
      RECT 3.755 1.815 3.945 2.875 ;
      RECT 4.94 0.83 5.13 2.875 ;
      RECT 3.755 2.685 5.13 2.875 ;
      RECT 9.41 0.425 10.395 0.62 ;
      RECT 6.615 1.55 6.805 1.83 ;
      RECT 10.085 0.425 10.275 1.83 ;
      RECT 6.615 1.64 10.275 1.83 ;
      RECT 9.63 1.64 9.82 2.265 ;
      RECT 7.68 1.64 7.87 2.285 ;
      RECT 11.46 2.26 13.16 2.45 ;
      RECT 11.015 0.43 12.95 0.62 ;
      RECT 12.76 0.955 14.385 1.145 ;
      RECT 12.76 0.43 12.95 1.99 ;
      RECT 10.91 1.8 12.95 1.99 ;
      RECT 10.91 1.8 11.1 2.45 ;
      RECT 10.555 2.26 11.1 2.45 ;
      RECT 14.1 0.43 14.775 0.62 ;
      RECT 13.35 1.79 16.125 1.98 ;
      RECT 14.585 0.43 14.775 2.475 ;
  END
END DSRNQV2_7TV50

MACRO FDCAP12_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FDCAP12_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.355 0.435 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 5.8 -0.12 6.08 0.635 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.575 0.52 0.78 1.92 ;
      RECT 5.275 1.07 5.465 2.48 ;
  END
END FDCAP12_7TV50

MACRO FDCAP4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FDCAP4_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.405 0.435 3.48 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.42 -0.12 1.7 0.565 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.565 0.365 0.765 2.045 ;
      RECT 1.05 1.065 1.28 1.345 ;
      RECT 1.05 1.065 1.24 2.48 ;
  END
END FDCAP4_7TV50

MACRO FDCAP8_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FDCAP8_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.395 0.435 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.885 -0.12 4.165 0.74 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.575 0.595 0.765 2.04 ;
      RECT 3.515 1.03 3.72 2.475 ;
  END
END FDCAP8_7TV50

MACRO FILLTIE_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLTIE_7TV50 0 0 ;
  SIZE 0.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.54 3.94 ;
      LAYER M1 ;
        RECT 0 3.24 0.96 3.48 ;
        RECT 0.38 2.33 0.57 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 0.26 1.46 ;
        RECT -0.12 -0.24 1.08 0.24 ;
        RECT 0.7 -0.24 1.08 1.46 ;
        RECT -0.12 1.08 1.08 1.46 ;
      LAYER M1 ;
        RECT 0 -0.12 0.96 0.12 ;
        RECT 0.335 -0.12 0.615 0.55 ;
    END
  END VSS
END FILLTIE_7TV50

MACRO F_DIODE2_7TV50
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN F_DIODE2_7TV50 0 0 ;
  SIZE 0.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.345 0.385 0.625 2.795 ;
        RECT 0.345 1.52 0.84 1.84 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 0.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 0.96 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.54 3.94 ;
    END
  END VNW
END F_DIODE2_7TV50

MACRO F_DIODEN2_7TV50
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN F_DIODEN2_7TV50 0 0 ;
  SIZE 0.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.32 0.32 0.84 1.29 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 0.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 0.96 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.54 3.94 ;
    END
  END VNW
END F_DIODEN2_7TV50

MACRO F_FILL16_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN F_FILL16_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.26 3.94 ;
    END
  END VNW
END F_FILL16_7TV50

MACRO F_FILL1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN F_FILL1_7TV50 0 0 ;
  SIZE 0.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 0.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 0.48 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 0.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.06 3.94 ;
    END
  END VNW
END F_FILL1_7TV50

MACRO F_FILL2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN F_FILL2_7TV50 0 0 ;
  SIZE 0.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 0.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 0.96 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 1.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.54 3.94 ;
    END
  END VNW
END F_FILL2_7TV50

MACRO F_FILL4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN F_FILL4_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
END F_FILL4_7TV50

MACRO F_FILL8_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN F_FILL8_7TV50 0 0 ;
  SIZE 3.84 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 3.24 3.84 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.12 3.84 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.96 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.42 3.94 ;
    END
  END VNW
END F_FILL8_7TV50

MACRO INV0P7_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV0P7_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.52 0.84 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.22 2.545 0.5 3.48 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.17 -0.12 0.45 0.765 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.115 0.595 1.305 2.475 ;
        RECT 1.08 1.52 1.32 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
END INV0P7_7TV50

MACRO INV16_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV16_7TV50 0 0 ;
  SIZE 15.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.28 1.56 7.6 1.8 ;
        RECT 7.165 1.61 9.395 1.8 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.855 2.4 1.135 3.48 ;
        RECT 2.555 2.79 2.835 3.48 ;
        RECT 4.255 2.79 4.535 3.48 ;
        RECT 5.995 2.79 6.275 3.48 ;
        RECT 7.735 2.79 8.015 3.48 ;
        RECT 9.49 2.79 9.77 3.48 ;
        RECT 11.19 2.79 11.47 3.48 ;
        RECT 12.89 2.79 13.17 3.48 ;
        RECT 14.59 2.395 14.87 3.48 ;
        RECT 0 3.24 15.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.305 -0.12 0.585 0.61 ;
        RECT 2.105 -0.12 2.385 0.565 ;
        RECT 3.905 -0.12 4.185 0.565 ;
        RECT 5.705 -0.12 5.985 0.565 ;
        RECT 7.505 -0.12 7.785 0.565 ;
        RECT 9.305 -0.12 9.585 0.565 ;
        RECT 11.105 -0.12 11.385 0.565 ;
        RECT 12.905 -0.12 13.185 0.565 ;
        RECT 14.75 -0.12 14.94 0.61 ;
        RECT 0 -0.12 15.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.25 0.595 1.44 0.955 ;
        RECT 3.05 0.595 3.24 0.955 ;
        RECT 4.85 0.595 5.04 0.955 ;
        RECT 6.65 0.595 6.84 0.955 ;
        RECT 8.45 0.595 8.64 0.955 ;
        RECT 10.225 0.765 10.415 2.475 ;
        RECT 10.25 0.595 10.44 0.955 ;
        RECT 10.16 1.56 10.49 1.8 ;
        RECT 12.05 0.595 12.24 0.955 ;
        RECT 1.705 2.285 14.02 2.475 ;
        RECT 13.85 0.595 14.04 0.955 ;
        RECT 1.25 0.765 14.04 0.955 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 15.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 15.94 3.94 ;
    END
  END VNW
END INV16_7TV50

MACRO INV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV1_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.12 1.04 0.36 1.36 ;
        RECT 0.12 1.17 0.835 1.36 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.23 2.36 0.51 3.48 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.18 -0.12 0.46 0.695 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.595 1.315 2.475 ;
        RECT 1.08 1.04 1.32 1.36 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
END INV1_7TV50

MACRO INV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV2_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.46 1.45 0.84 1.865 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.32 0.485 3.48 ;
        RECT 1.955 2.3 2.235 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.61 ;
        RECT 1.955 -0.12 2.235 0.61 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.56 1.29 2.475 ;
        RECT 1.08 0.56 1.32 0.88 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
END INV2_7TV50

MACRO INV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV3_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.785 1.56 1.365 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.4 0.435 3.48 ;
        RECT 2.005 2.795 2.285 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.61 ;
        RECT 1.955 -0.12 2.235 0.565 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.595 1.29 0.955 ;
        RECT 2 0.765 2.19 2.43 ;
        RECT 2 1.56 2.33 1.8 ;
        RECT 2.9 0.595 3.09 0.955 ;
        RECT 1.1 0.765 3.09 0.955 ;
        RECT 1.005 2.24 3.135 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
END INV3_7TV50

MACRO INV4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV4_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.53 1.56 1.155 1.84 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.305 2.405 0.585 3.48 ;
        RECT 2.005 2.795 2.285 3.48 ;
        RECT 3.755 2.405 4.035 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.565 ;
        RECT 1.955 -0.12 2.235 0.565 ;
        RECT 3.755 -0.12 4.035 0.565 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.595 1.29 0.955 ;
        RECT 2.07 0.765 2.26 2.43 ;
        RECT 2 1.56 2.33 1.8 ;
        RECT 2.9 0.595 3.09 0.955 ;
        RECT 1.1 0.765 3.09 0.955 ;
        RECT 1.155 2.24 3.135 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
END INV4_7TV50

MACRO INV6_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV6_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.56 2.91 1.8 ;
        RECT 2.24 1.61 2.91 1.8 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.455 2.355 0.735 3.48 ;
        RECT 2.155 2.79 2.435 3.48 ;
        RECT 3.855 2.79 4.135 3.48 ;
        RECT 5.575 2.34 5.855 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.175 -0.12 0.455 0.61 ;
        RECT 1.975 -0.12 2.255 0.565 ;
        RECT 3.775 -0.12 4.055 0.565 ;
        RECT 5.575 -0.12 5.855 0.61 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.12 0.56 1.31 0.955 ;
        RECT 2.92 0.595 3.11 0.955 ;
        RECT 3.44 0.765 3.63 2.49 ;
        RECT 3.44 1.56 3.77 1.8 ;
        RECT 4.72 0.595 4.91 0.955 ;
        RECT 1.12 0.765 4.91 0.955 ;
        RECT 1.305 2.3 4.985 2.49 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
END INV6_7TV50

MACRO INV8_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV8_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.92 1.56 4.24 1.8 ;
        RECT 3.64 1.61 4.7 1.8 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.7 2.35 0.98 3.48 ;
        RECT 2.4 2.795 2.68 3.48 ;
        RECT 4.115 2.795 4.395 3.48 ;
        RECT 5.815 2.795 6.095 3.48 ;
        RECT 7.515 2.35 7.795 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.315 -0.12 0.595 0.61 ;
        RECT 2.115 -0.12 2.395 0.565 ;
        RECT 3.915 -0.12 4.195 0.565 ;
        RECT 5.715 -0.12 5.995 0.565 ;
        RECT 7.515 -0.12 7.795 0.61 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.595 1.45 0.955 ;
        RECT 3.06 0.595 3.25 0.955 ;
        RECT 4.86 0.595 5.05 0.955 ;
        RECT 5.36 1.56 5.69 1.8 ;
        RECT 5.5 0.765 5.69 2.55 ;
        RECT 6.66 0.595 6.85 0.955 ;
        RECT 1.26 0.765 6.85 0.955 ;
        RECT 1.55 2.36 6.945 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
END INV8_7TV50

MACRO LAHQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LAHQV1_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.92 1.56 3.52 1.8 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.915 1.5 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.28 1.52 8.57 1.84 ;
        RECT 8.38 0.595 8.57 2.5 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.745 1.345 3.48 ;
        RECT 2.82 2.52 3.055 3.48 ;
        RECT 6.035 2.28 6.315 3.48 ;
        RECT 7.485 2.28 7.765 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 2.545 -0.12 2.825 0.875 ;
        RECT 5.945 -0.12 6.225 0.875 ;
        RECT 7.435 -0.12 7.715 0.875 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 4.005 1.76 4.195 2.32 ;
      RECT 2.41 2.13 4.195 2.32 ;
      RECT 0.2 2.285 1.735 2.475 ;
      RECT 1.545 1.76 1.735 2.865 ;
      RECT 2.41 2.13 2.6 2.865 ;
      RECT 1.545 2.675 2.6 2.865 ;
      RECT 1.955 0.625 2.235 0.815 ;
      RECT 2.02 1.075 5.045 1.265 ;
      RECT 4.855 1.075 5.045 2.04 ;
      RECT 2.02 0.625 2.21 2.475 ;
      RECT 4.245 0.64 5.435 0.83 ;
      RECT 5.245 1.075 6.48 1.265 ;
      RECT 5.245 0.64 5.435 2.43 ;
      RECT 4.435 2.24 5.435 2.43 ;
      RECT 6.535 0.64 6.87 0.83 ;
      RECT 5.66 1.745 6.87 1.935 ;
      RECT 6.68 0.64 6.87 2.475 ;
  END
END LAHQV1_7TV50

MACRO LAHQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LAHQV2_7TV50 0 0 ;
  SIZE 10.08 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.92 1.56 3.52 1.8 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.915 1.5 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.28 1.52 8.57 1.84 ;
        RECT 8.38 0.595 8.57 2.5 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.745 1.345 3.48 ;
        RECT 2.82 2.685 3.055 3.48 ;
        RECT 6.035 2.28 6.315 3.48 ;
        RECT 7.485 2.28 7.765 3.48 ;
        RECT 9.185 2.22 9.465 3.48 ;
        RECT 0 3.24 10.08 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 2.545 -0.12 2.825 0.79 ;
        RECT 5.945 -0.12 6.225 0.875 ;
        RECT 7.435 -0.12 7.715 0.875 ;
        RECT 9.235 -0.12 9.515 0.75 ;
        RECT 0 -0.12 10.08 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 10.2 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 10.66 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 4.005 1.76 4.195 2.32 ;
      RECT 2.41 2.13 4.195 2.32 ;
      RECT 0.2 2.285 1.735 2.475 ;
      RECT 1.545 1.76 1.735 2.865 ;
      RECT 2.41 2.13 2.6 2.865 ;
      RECT 1.545 2.675 2.6 2.865 ;
      RECT 1.955 0.64 2.235 0.83 ;
      RECT 2.02 1.075 5.045 1.265 ;
      RECT 4.855 1.075 5.045 2.04 ;
      RECT 2.02 0.64 2.21 2.475 ;
      RECT 4.245 0.64 5.435 0.83 ;
      RECT 5.245 1.075 6.48 1.265 ;
      RECT 5.245 0.64 5.435 2.43 ;
      RECT 4.435 2.24 5.435 2.43 ;
      RECT 6.535 0.64 6.87 0.83 ;
      RECT 5.66 1.745 6.87 1.935 ;
      RECT 6.68 0.64 6.87 2.475 ;
  END
END LAHQV2_7TV50

MACRO LAHRNQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LAHRNQV1_7TV50 0 0 ;
  SIZE 10.56 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.38 1.905 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.91 1.505 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.13 0.56 10.32 2.475 ;
        RECT 10.13 0.56 10.44 0.88 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.11 2 7.56 2.32 ;
    END
  END RDN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.285 1.285 3.48 ;
        RECT 3.425 2.38 3.705 3.48 ;
        RECT 6.745 2.97 7.025 3.48 ;
        RECT 9.235 2.275 9.515 3.48 ;
        RECT 0 3.24 10.56 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 6.835 -0.12 7.115 0.695 ;
        RECT 9.225 -0.12 9.505 0.875 ;
        RECT 0 -0.12 10.56 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.27 -0.24 4.86 1.53 ;
        RECT -0.12 -0.24 10.68 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.27 3.94 ;
        RECT 4.86 1.46 11.14 3.94 ;
        RECT -0.58 1.53 11.14 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.775 1.66 1.965 ;
      RECT 0.2 0.595 0.39 2.48 ;
      RECT 2 0.595 2.19 1.335 ;
      RECT 1.9 1.145 4.115 1.335 ;
      RECT 1.9 1.145 2.09 2.54 ;
      RECT 4.795 0.895 4.985 2.07 ;
      RECT 4.705 1.88 4.985 2.07 ;
      RECT 2.665 0.32 6.265 0.51 ;
      RECT 6.075 0.32 6.265 1.085 ;
      RECT 2.665 0.32 2.855 0.9 ;
      RECT 2.575 0.71 2.855 0.9 ;
      RECT 7.78 0.46 7.97 1.085 ;
      RECT 6.075 0.895 7.97 1.085 ;
      RECT 6.31 1.445 8.56 1.635 ;
      RECT 8.37 0.595 8.56 2.475 ;
      RECT 4.275 0.71 4.555 0.9 ;
      RECT 4.315 0.71 4.505 2.77 ;
      RECT 4.315 2.58 7.89 2.77 ;
      RECT 7.7 2.755 8.98 2.945 ;
  END
END LAHRNQV1_7TV50

MACRO LAHRNQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LAHRNQV2_7TV50 0 0 ;
  SIZE 11.52 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.38 1.905 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.91 1.505 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.13 0.56 10.32 2.475 ;
        RECT 10.13 0.56 10.44 0.88 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.11 2 7.56 2.32 ;
    END
  END RDN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.285 1.285 3.48 ;
        RECT 3.425 2.38 3.705 3.48 ;
        RECT 6.745 2.97 7.025 3.48 ;
        RECT 9.235 2.275 9.515 3.48 ;
        RECT 10.995 2.275 11.275 3.48 ;
        RECT 0 3.24 11.52 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 6.835 -0.12 7.115 0.695 ;
        RECT 9.225 -0.12 9.505 0.875 ;
        RECT 11.025 -0.12 11.305 0.785 ;
        RECT 0 -0.12 11.52 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.27 -0.24 4.86 1.53 ;
        RECT -0.12 -0.24 11.64 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.27 3.94 ;
        RECT 4.86 1.46 12.1 3.94 ;
        RECT -0.58 1.53 12.1 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.775 1.66 1.965 ;
      RECT 0.2 0.595 0.39 2.48 ;
      RECT 2 0.595 2.19 1.335 ;
      RECT 1.9 1.145 4.115 1.335 ;
      RECT 1.9 1.145 2.09 2.54 ;
      RECT 4.795 0.895 4.985 2.07 ;
      RECT 4.705 1.88 4.985 2.07 ;
      RECT 2.665 0.32 6.265 0.51 ;
      RECT 6.075 0.32 6.265 1.085 ;
      RECT 2.665 0.32 2.855 0.9 ;
      RECT 2.575 0.71 2.855 0.9 ;
      RECT 7.78 0.46 7.97 1.085 ;
      RECT 6.075 0.895 7.97 1.085 ;
      RECT 6.31 1.445 8.56 1.635 ;
      RECT 8.37 0.595 8.56 2.475 ;
      RECT 4.275 0.71 4.555 0.9 ;
      RECT 4.315 0.71 4.505 2.77 ;
      RECT 4.315 2.58 7.89 2.77 ;
      RECT 7.7 2.695 8.98 2.885 ;
  END
END LAHRNQV2_7TV50

MACRO LAHSQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LAHSQV1_7TV50 0 0 ;
  SIZE 10.08 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.92 1.56 3.28 1.96 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.59 1.04 1.04 1.36 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.28 0.6 9.47 2.48 ;
        RECT 9.2 0.6 9.52 0.84 ;
    END
  END Q
  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.025 1.89 7.285 2.28 ;
        RECT 6.8 2.04 7.285 2.28 ;
    END
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.22 1.285 3.48 ;
        RECT 6.765 2.75 7.045 3.48 ;
        RECT 8.385 2.28 8.665 3.48 ;
        RECT 0 3.24 10.08 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.81 ;
        RECT 2.545 -0.12 2.825 0.73 ;
        RECT 5.945 -0.12 6.225 0.685 ;
        RECT 8.335 -0.12 8.615 0.67 ;
        RECT 0 -0.12 10.08 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.405 1.46 ;
        RECT -0.12 -0.24 10.2 1.315 ;
        RECT 7.36 -0.24 10.2 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 5.405 1.315 7.36 3.94 ;
        RECT -0.58 1.46 10.66 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.76 1.66 1.95 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 2 0.595 2.19 1.12 ;
      RECT 1.9 0.93 4 1.12 ;
      RECT 1.9 0.93 2.09 2.475 ;
      RECT 4.665 0.885 4.855 2.07 ;
      RECT 3.725 1.88 4.855 2.07 ;
      RECT 2.49 2.38 2.68 2.895 ;
      RECT 5.915 2.07 6.105 2.895 ;
      RECT 2.49 2.705 6.105 2.895 ;
      RECT 4.245 0.495 5.33 0.685 ;
      RECT 6.89 0.45 7.08 1.12 ;
      RECT 5.14 0.93 7.37 1.12 ;
      RECT 5.14 0.495 5.33 2.505 ;
      RECT 4.1 2.315 5.33 2.505 ;
      RECT 7.435 0.495 7.77 0.685 ;
      RECT 7.57 0.495 7.77 1.62 ;
      RECT 5.57 1.43 7.77 1.62 ;
      RECT 7.58 0.495 7.77 2.48 ;
  END
END LAHSQV1_7TV50

MACRO LAHSQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LAHSQV2_7TV50 0 0 ;
  SIZE 11.04 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.92 1.56 3.28 1.96 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.59 1.04 1.04 1.36 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.6 0.525 9.79 2.48 ;
        RECT 9.6 0.525 9.96 0.88 ;
    END
  END Q
  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.095 1.86 7.285 2.28 ;
        RECT 6.8 2.04 7.285 2.28 ;
    END
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.22 1.285 3.48 ;
        RECT 6.765 2.75 7.045 3.48 ;
        RECT 8.705 2.28 8.985 3.48 ;
        RECT 10.405 2.31 10.685 3.48 ;
        RECT 0 3.24 11.04 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.83 ;
        RECT 2.545 -0.12 2.825 0.7 ;
        RECT 5.945 -0.12 6.225 0.655 ;
        RECT 8.655 -0.12 8.935 0.705 ;
        RECT 10.455 -0.12 10.735 0.705 ;
        RECT 0 -0.12 11.04 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.37 1.46 ;
        RECT -0.12 -0.24 11.16 1.285 ;
        RECT 7.395 -0.24 11.16 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 5.37 1.285 7.395 3.94 ;
        RECT -0.58 1.46 11.62 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.805 1.66 1.995 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 2 0.595 2.19 1.12 ;
      RECT 1.9 0.93 4 1.12 ;
      RECT 1.9 0.93 2.09 2.475 ;
      RECT 4.665 0.855 4.855 2.07 ;
      RECT 3.725 1.88 4.855 2.07 ;
      RECT 2.49 2.38 2.68 2.895 ;
      RECT 5.915 2.04 6.105 2.895 ;
      RECT 2.49 2.705 6.105 2.895 ;
      RECT 4.245 0.465 5.33 0.655 ;
      RECT 6.89 0.42 7.08 1.195 ;
      RECT 5.14 1.005 7.69 1.195 ;
      RECT 5.14 0.465 5.33 2.505 ;
      RECT 4.1 2.315 5.33 2.505 ;
      RECT 7.755 0.57 8.09 0.76 ;
      RECT 7.89 0.57 8.09 1.64 ;
      RECT 5.57 1.45 8.09 1.64 ;
      RECT 7.9 0.57 8.09 2.48 ;
  END
END LAHSQV2_7TV50

MACRO MAJ23V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJ23V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.04 0.925 1.32 ;
        RECT 0.56 1.04 3.63 1.23 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.695 1.825 1.885 2.19 ;
        RECT 1.695 2 2.76 2.19 ;
        RECT 2.57 2 2.76 2.97 ;
        RECT 2.52 2.48 2.76 2.8 ;
        RECT 4.22 1.825 4.41 2.97 ;
        RECT 2.57 2.78 4.41 2.97 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.465 2.935 1.8 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 2.9 1.395 3.48 ;
        RECT 4.61 2.42 4.845 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 -0.12 1.395 0.45 ;
        RECT 4.675 -0.12 4.955 0.76 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.62 0.525 5.81 2.44 ;
        RECT 5.4 2 5.81 2.44 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.205 2.435 2.305 2.625 ;
      RECT 0.155 0.57 0.435 0.84 ;
      RECT 2.075 0.57 2.355 0.84 ;
      RECT 0.155 0.65 2.355 0.84 ;
      RECT 2.975 0.57 4.02 0.76 ;
      RECT 3.83 1.005 5.22 1.195 ;
      RECT 3.83 0.57 4.02 2.525 ;
      RECT 2.96 2.335 4.02 2.525 ;
  END
END MAJ23V1_7TV50

MACRO MAJ23V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJ23V2_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.04 0.88 1.32 ;
        RECT 0.56 1.04 3.48 1.23 ;
        RECT 3.2 1.04 3.48 1.27 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.745 1.905 1.935 2.19 ;
        RECT 1.745 2 2.7 2.19 ;
        RECT 2.51 2 2.7 2.97 ;
        RECT 2.51 2.48 2.76 2.97 ;
        RECT 4.22 1.815 4.41 2.97 ;
        RECT 2.51 2.78 4.41 2.97 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.43 2.87 1.8 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.165 2.795 1.445 3.48 ;
        RECT 4.67 2.75 4.93 3.48 ;
        RECT 6.325 2.405 6.605 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 -0.12 1.395 0.45 ;
        RECT 4.675 -0.12 4.955 0.565 ;
        RECT 6.475 -0.12 6.755 0.565 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 2 5.815 2.32 ;
        RECT 5.62 0.525 5.815 2.48 ;
        RECT 5.52 2 5.815 2.48 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.205 2.39 2.31 2.58 ;
      RECT 2.12 2.39 2.31 2.67 ;
      RECT 0.155 0.47 0.435 0.84 ;
      RECT 2.075 0.47 2.355 0.84 ;
      RECT 0.155 0.65 2.355 0.84 ;
      RECT 2.975 0.505 3.96 0.695 ;
      RECT 3.77 1.225 5.15 1.415 ;
      RECT 3.77 0.505 3.96 2.495 ;
      RECT 3.025 2.305 3.96 2.495 ;
  END
END MAJ23V2_7TV50

MACRO MAOI222V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAOI222V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.395 1.56 4.745 1.8 ;
        RECT 3.78 1.56 4.91 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.08 1.84 1.32 ;
        RECT 1.48 1.13 5.66 1.32 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.56 2.83 1.8 ;
        RECT 0.63 1.56 3.11 1.75 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.355 0.435 3.48 ;
        RECT 1.855 2.745 2.135 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.685 ;
        RECT 2.445 -0.12 2.725 0.435 ;
        RECT 5.965 -0.12 6.245 0.435 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.855 0.64 6.12 0.83 ;
        RECT 5.88 0.64 6.12 2.43 ;
        RECT 5.105 2.24 6.12 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.24 3.585 2.43 ;
      RECT 2.455 2.75 6.235 2.94 ;
  END
END MAOI222V1_7TV50

MACRO MAOI222V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAOI222V2_7TV50 0 0 ;
  SIZE 11.52 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.255 1.415 7.805 1.605 ;
        RECT 7.615 1.415 7.805 1.85 ;
        RECT 8.72 1.56 9.04 1.85 ;
        RECT 7.615 1.66 9.955 1.85 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.075 1.84 1.32 ;
        RECT 1.48 1.13 4.77 1.32 ;
        RECT 4.58 1.025 8.22 1.215 ;
        RECT 8.03 1.075 10.48 1.265 ;
        RECT 10.29 1.075 10.48 1.63 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.92 1.56 4.27 1.995 ;
        RECT 0.63 1.805 7.41 1.995 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.355 0.435 3.48 ;
        RECT 1.855 2.745 2.135 3.48 ;
        RECT 3.555 2.745 3.835 3.48 ;
        RECT 0 3.24 11.52 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.685 ;
        RECT 3.72 -0.12 4 0.39 ;
        RECT 7.565 -0.12 7.845 0.39 ;
        RECT 11.085 -0.12 11.365 0.39 ;
        RECT 0 -0.12 11.52 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.855 0.59 10.92 0.78 ;
        RECT 10.68 0.59 10.92 2.43 ;
        RECT 8.455 2.24 10.92 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 11.64 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 12.1 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.005 2.355 7.035 2.545 ;
      RECT 4.205 2.75 11.285 2.94 ;
  END
END MAOI222V2_7TV50

MACRO MOAI222V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MOAI222V1_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.875 2.32 2.28 ;
        RECT 1.825 1.875 2.855 2.065 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.23 1.32 1.84 ;
        RECT 1.08 1.23 5.375 1.42 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.84 1.56 6.175 1.81 ;
        RECT 3.625 1.62 6.175 1.81 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 2.595 0.4 3.48 ;
        RECT 3.92 2.97 4.2 3.48 ;
        RECT 6.37 2.355 6.65 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.66 -0.12 4.94 0.435 ;
        RECT 6.52 -0.12 6.8 0.685 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.65 0.84 0.84 2.67 ;
        RECT 1.19 0.71 1.47 1.03 ;
        RECT 0.65 0.84 1.47 1.03 ;
        RECT 0.65 2.48 5.05 2.67 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.605 -0.24 3.975 1.53 ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.605 3.94 ;
        RECT 3.975 1.46 7.78 3.94 ;
        RECT -0.58 1.53 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.23 0.32 4.35 0.51 ;
      RECT 0.23 0.32 0.51 0.64 ;
      RECT 2.15 0.32 2.43 0.64 ;
      RECT 4.07 0.32 4.35 0.64 ;
      RECT 3.11 0.71 3.39 1.03 ;
      RECT 5.665 0.595 5.855 1.03 ;
      RECT 3.11 0.84 5.855 1.03 ;
  END
END MOAI222V1_7TV50

MACRO MOAI222V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MOAI222V2_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.875 2.32 2.28 ;
        RECT 1.75 1.875 4.16 2.065 ;
        RECT 3.97 1.99 6.64 2.18 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.21 1.32 1.84 ;
        RECT 1.08 1.21 10.9 1.4 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.12 1.56 11.44 1.8 ;
        RECT 4.46 1.6 11.64 1.79 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.455 2.91 0.735 3.48 ;
        RECT 3.805 2.845 4.085 3.48 ;
        RECT 7.77 2.845 8.05 3.48 ;
        RECT 8.385 2.845 8.665 3.48 ;
        RECT 12.045 2.245 12.325 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 8.445 -0.12 8.725 0.62 ;
        RECT 10.245 -0.12 10.525 0.62 ;
        RECT 12.045 -0.12 12.325 0.665 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.65 0.82 0.84 2.71 ;
        RECT 1.135 0.71 1.415 1.01 ;
        RECT 0.65 2.52 2.695 2.71 ;
        RECT 3.055 0.71 3.335 1.01 ;
        RECT 0.65 0.82 3.335 1.01 ;
        RECT 5.81 2.455 6.09 2.845 ;
        RECT 2.505 2.455 10.47 2.645 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.58 -0.24 7.68 1.53 ;
        RECT -0.12 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.58 3.94 ;
        RECT 7.68 1.46 13.06 3.94 ;
        RECT -0.58 1.53 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.175 0.32 8.135 0.51 ;
      RECT 0.175 0.32 0.455 0.62 ;
      RECT 2.095 0.32 2.375 0.62 ;
      RECT 4.015 0.32 4.295 0.62 ;
      RECT 5.935 0.32 6.215 0.62 ;
      RECT 7.855 0.32 8.135 0.62 ;
      RECT 4.975 0.71 5.255 1.01 ;
      RECT 6.895 0.71 7.175 1.01 ;
      RECT 9.39 0.58 9.58 1.01 ;
      RECT 11.19 0.58 11.38 1.01 ;
      RECT 4.975 0.82 11.38 1.01 ;
  END
END MOAI222V2_7TV50

MACRO MUX2NV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2NV1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.515 0.9 1.995 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.56 1.8 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.395 1.075 4.24 1.265 ;
        RECT 3.92 1.075 4.24 1.32 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.22 2.24 0.5 3.48 ;
        RECT 3.42 2.4 3.7 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.17 -0.12 0.455 0.735 ;
        RECT 3.57 -0.12 3.85 0.875 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.865 0.56 2.055 2.475 ;
        RECT 1.865 0.56 2.28 0.88 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.255 1.76 2.445 2.19 ;
      RECT 4.515 0.595 4.705 2.19 ;
      RECT 2.255 2 4.705 2.19 ;
      RECT 4.315 2 4.505 2.475 ;
  END
END MUX2NV1_7TV50

MACRO MUX2NV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2NV2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 1.515 0.895 1.84 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.315 1.56 6.915 1.8 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.415 5.745 1.84 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.04 2.725 1.32 3.48 ;
        RECT 4.18 2.97 4.46 3.48 ;
        RECT 5.985 2.69 6.22 3.48 ;
        RECT 7.64 2.275 7.92 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.34 -0.12 1.62 0.625 ;
        RECT 5.59 -0.12 5.87 0.565 ;
        RECT 7.39 -0.12 7.67 0.71 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.785 1.56 2.975 2.57 ;
        RECT 3.2 0.735 3.39 1.8 ;
        RECT 2.785 1.56 3.39 1.8 ;
        RECT 3.2 0.735 3.48 0.925 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.855 -0.24 4.73 1.555 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.855 3.94 ;
        RECT 4.73 1.46 8.74 3.94 ;
        RECT -0.58 1.555 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.235 2.335 2.17 2.525 ;
      RECT 0.235 2.335 0.425 3.03 ;
      RECT 0.485 0.595 0.675 1.015 ;
      RECT 2.285 0.595 2.475 1.015 ;
      RECT 0.485 0.825 2.475 1.015 ;
      RECT 2.81 0.32 4.97 0.51 ;
      RECT 4.69 0.32 4.97 0.565 ;
      RECT 2.81 0.32 3 1.31 ;
      RECT 3.69 0.32 3.88 2.205 ;
      RECT 3.69 2.015 5.28 2.205 ;
      RECT 5.09 2.015 5.28 2.65 ;
      RECT 5.09 2.46 5.37 2.65 ;
      RECT 4.1 0.735 4.38 0.955 ;
      RECT 6.535 0.53 6.725 0.955 ;
      RECT 4.1 0.765 6.725 0.955 ;
      RECT 5.57 2.3 7.07 2.49 ;
      RECT 3.59 2.58 4.885 2.77 ;
      RECT 4.695 2.58 4.885 3.04 ;
      RECT 5.57 2.3 5.76 3.04 ;
      RECT 4.695 2.85 5.76 3.04 ;
  END
END MUX2NV2_7TV50

MACRO MUX2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.08 1.08 4.72 1.32 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.52 1.8 1.97 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.91 1.985 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.24 1.285 3.48 ;
        RECT 4.265 2.275 4.545 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 4.455 -0.12 4.735 0.875 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.16 0.56 5.35 2.475 ;
        RECT 5.16 0.56 5.64 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.075 3.45 1.265 ;
      RECT 2.175 1.075 2.365 2.04 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 2.755 0.64 3.84 0.83 ;
      RECT 3.65 0.64 3.84 1.995 ;
      RECT 2.65 1.805 4.92 1.995 ;
      RECT 2.65 1.805 2.84 2.475 ;
  END
END MUX2V1_7TV50

MACRO MUX2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2V2_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.08 1.08 4.72 1.32 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 1.56 1.84 1.8 ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.6 1.075 2.51 1.265 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.425 1.285 3.48 ;
        RECT 4.265 2.275 4.545 3.48 ;
        RECT 5.965 2.275 6.245 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 4.455 -0.12 4.735 0.745 ;
        RECT 6.255 -0.12 6.535 0.75 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.16 0.56 5.35 2.475 ;
        RECT 5.16 0.56 5.64 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.215 1.03 3.405 1.945 ;
      RECT 2.175 1.755 3.405 1.945 ;
      RECT 2.175 1.755 2.365 2.19 ;
      RECT 0.2 2 2.365 2.19 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 2.755 0.64 3.84 0.83 ;
      RECT 3.65 1.805 4.92 1.995 ;
      RECT 3.65 0.64 3.84 2.43 ;
      RECT 2.605 2.24 3.84 2.43 ;
  END
END MUX2V2_7TV50

MACRO MUX3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX3V1_7TV50 0 0 ;
  SIZE 10.08 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.08 1.08 4.72 1.32 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.435 1.56 1.84 1.92 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.18 1.03 8.62 1.36 ;
    END
  END I2
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.88 2.04 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.38 1.08 6.57 2.255 ;
        RECT 6.38 1.08 7.12 1.32 ;
        RECT 6.38 1.08 7.5 1.27 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.245 1.285 3.48 ;
        RECT 4.265 2.275 4.5 3.48 ;
        RECT 8.45 2.42 8.73 3.48 ;
        RECT 0 3.24 10.08 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 4.455 -0.12 4.735 0.865 ;
        RECT 8.545 -0.12 8.825 0.82 ;
        RECT 0 -0.12 10.08 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.345 0.6 9.535 2.475 ;
        RECT 9.2 0.6 9.725 0.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 10.2 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 10.66 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.075 3.45 1.265 ;
      RECT 2.175 1.075 2.365 2.055 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.4 1.03 5.785 1.31 ;
      RECT 5.4 0.595 5.59 2.43 ;
      RECT 5.115 2.24 5.59 2.43 ;
      RECT 2.755 0.64 3.84 0.83 ;
      RECT 3.65 1.805 4.89 1.995 ;
      RECT 3.65 0.64 3.84 2.43 ;
      RECT 2.605 2.24 3.84 2.43 ;
      RECT 4.7 1.805 4.89 2.82 ;
      RECT 5.99 0.595 6.18 2.82 ;
      RECT 4.7 2.63 6.18 2.82 ;
      RECT 6.845 0.64 7.91 0.83 ;
      RECT 7.72 1.805 9.105 1.995 ;
      RECT 7.72 0.64 7.91 2.645 ;
      RECT 6.795 2.455 7.91 2.645 ;
  END
END MUX3V1_7TV50

MACRO MUX3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX3V2_7TV50 0 0 ;
  SIZE 11.04 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.08 1.08 4.72 1.32 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.52 1.8 1.97 ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.18 1.03 8.62 1.36 ;
    END
  END I2
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.91 1.985 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.38 1.08 6.57 2.255 ;
        RECT 6.38 1.08 7.12 1.32 ;
        RECT 6.38 1.08 7.5 1.27 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.245 1.285 3.48 ;
        RECT 4.265 2.275 4.5 3.48 ;
        RECT 8.45 2.375 8.73 3.48 ;
        RECT 10.15 2.275 10.43 3.48 ;
        RECT 0 3.24 11.04 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 4.455 -0.12 4.735 0.865 ;
        RECT 8.545 -0.12 8.825 0.82 ;
        RECT 10.345 -0.12 10.625 0.75 ;
        RECT 0 -0.12 11.04 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.345 0.6 9.535 2.475 ;
        RECT 9.2 0.6 9.725 0.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 11.16 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 11.62 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.075 3.45 1.265 ;
      RECT 2.175 1.075 2.365 2.055 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.4 1.03 5.785 1.31 ;
      RECT 5.4 0.595 5.59 2.43 ;
      RECT 5.115 2.24 5.59 2.43 ;
      RECT 2.755 0.64 3.84 0.83 ;
      RECT 3.65 1.805 4.89 1.995 ;
      RECT 3.65 0.64 3.84 2.43 ;
      RECT 2.605 2.24 3.84 2.43 ;
      RECT 4.7 1.805 4.89 2.82 ;
      RECT 5.99 0.595 6.18 2.82 ;
      RECT 4.7 2.63 6.18 2.82 ;
      RECT 6.845 0.64 7.91 0.83 ;
      RECT 7.72 1.805 9.105 1.995 ;
      RECT 7.72 0.64 7.91 2.69 ;
      RECT 6.795 2.5 7.91 2.69 ;
  END
END MUX3V2_7TV50

MACRO NAND2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2V1_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 2.005 1.875 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.315 1.52 0.84 1.84 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.75 0.485 3.48 ;
        RECT 1.915 2.75 2.195 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.61 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.56 1.29 2.475 ;
        RECT 1.08 0.56 1.32 0.88 ;
        RECT 1.08 0.56 2.195 0.75 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
END NAND2V1_7TV50

MACRO NAND2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.425 1.08 2.005 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.56 2.8 1.8 ;
        RECT 0.63 1.61 3.28 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.75 0.435 3.48 ;
        RECT 1.905 2.795 2.185 3.48 ;
        RECT 3.655 2.795 3.935 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 -0.12 0.485 0.61 ;
        RECT 3.605 -0.12 3.885 0.565 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.905 0.64 3 0.83 ;
        RECT 2.81 0.83 3.8 1.02 ;
        RECT 3.48 0.83 3.8 1.36 ;
        RECT 3.61 0.83 3.8 2.435 ;
        RECT 1.005 2.245 3.8 2.435 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
END NAND2V2_7TV50

MACRO NAND2V3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2V3_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.08 3.28 1.32 ;
        RECT 2.41 1.13 5.41 1.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.94 1.56 1.49 1.8 ;
        RECT 0.94 1.61 3.415 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.36 0.565 3.48 ;
        RECT 2.025 2.795 2.305 3.48 ;
        RECT 3.84 2.795 4.12 3.48 ;
        RECT 5.605 2.795 5.885 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.335 -0.12 0.615 0.61 ;
        RECT 3.795 -0.12 4.075 0.39 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 0.6 3.76 0.84 ;
        RECT 2.035 0.6 5.885 0.79 ;
        RECT 5.695 0.6 5.885 2.435 ;
        RECT 1.135 2.245 5.885 2.435 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
END NAND2V3_7TV50

MACRO NAND2V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2V4_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.08 2.8 1.32 ;
        RECT 2.09 1.08 5.145 1.27 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.92 1.56 4.24 1.8 ;
        RECT 0.65 1.61 6.945 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.22 2.75 0.5 3.48 ;
        RECT 1.92 2.795 2.2 3.48 ;
        RECT 3.67 2.795 3.95 3.48 ;
        RECT 5.44 2.795 5.72 3.48 ;
        RECT 7.14 2.795 7.42 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.61 ;
        RECT 3.62 -0.12 3.91 0.39 ;
        RECT 7.15 -0.12 7.43 0.39 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 0.6 3.76 0.84 ;
        RECT 1.87 0.6 7.34 0.79 ;
        RECT 7.145 0.6 7.34 2.445 ;
        RECT 1.07 2.255 7.34 2.445 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.26 3.94 ;
    END
  END VNW
END NAND2V4_7TV50

MACRO NAND2XBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2XBV1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.03 2.5 1.36 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.525 1.52 0.84 1.98 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.4 0.435 3.48 ;
        RECT 1.855 2.42 2.135 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.965 -0.12 2.245 0.39 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.205 0.64 1.24 0.83 ;
        RECT 0.56 0.6 0.88 0.84 ;
        RECT 0.56 0.64 1.24 0.84 ;
        RECT 1.05 0.64 1.24 2.475 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.575 1.005 1.765 1.92 ;
      RECT 2.97 0.595 3.16 1.92 ;
      RECT 1.575 1.73 3.16 1.92 ;
      RECT 2.75 1.73 2.94 2.475 ;
  END
END NAND2XBV1_7TV50

MACRO NAND2XBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2XBV2_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.925 1.475 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.2 1.08 2.8 1.36 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.09 2.36 1.37 3.48 ;
        RECT 2.91 2.785 3.19 3.48 ;
        RECT 4.66 2.795 4.94 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.15 -0.12 1.43 0.39 ;
        RECT 4.61 -0.12 4.89 0.595 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.955 0.595 3.41 0.875 ;
        RECT 3.22 0.795 4.825 0.985 ;
        RECT 4.635 0.795 4.825 2.43 ;
        RECT 2.06 2.24 4.825 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.19 0.64 1.97 0.83 ;
      RECT 1.78 0.64 1.97 1.75 ;
      RECT 4.245 1.47 4.435 1.75 ;
      RECT 1.78 1.56 4.435 1.75 ;
      RECT 0.19 0.64 0.39 2.43 ;
      RECT 0.19 2.24 0.52 2.43 ;
  END
END NAND2XBV2_7TV50

MACRO NAND2XBV4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2XBV4_7TV50 0 0 ;
  SIZE 9.6 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.84 2.04 ;
        RECT 0.6 1.76 0.96 2.04 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.03 3.24 1.605 ;
        RECT 3 1.415 7.115 1.605 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.51 2.545 0.79 3.48 ;
        RECT 2.21 2.545 2.49 3.48 ;
        RECT 3.91 2.765 4.19 3.48 ;
        RECT 5.61 2.765 5.89 3.48 ;
        RECT 7.31 2.765 7.59 3.48 ;
        RECT 9.01 2.755 9.29 3.48 ;
        RECT 0 3.24 9.6 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.24 -0.12 0.52 0.83 ;
        RECT 2.1 -0.12 2.38 0.83 ;
        RECT 5.56 -0.12 5.84 0.63 ;
        RECT 9.02 -0.12 9.3 0.63 ;
        RECT 0 -0.12 9.6 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.905 0.595 4.095 1.205 ;
        RECT 7.305 0.595 7.495 1.205 ;
        RECT 3.905 1.015 9.205 1.205 ;
        RECT 8.72 1.015 9.205 1.32 ;
        RECT 9.015 1.015 9.205 2.55 ;
        RECT 3.06 2.36 9.205 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 9.72 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 10.18 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.185 0.595 1.375 1.995 ;
      RECT 1.185 1.805 8.815 1.995 ;
      RECT 1.405 1.805 1.595 2.535 ;
  END
END NAND2XBV4_7TV50

MACRO NAND3BBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBV1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.755 1.56 5.2 1.885 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.93 1.965 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.53 1.52 1.86 1.965 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.12 2.42 1.4 3.48 ;
        RECT 2.89 2.79 3.17 3.48 ;
        RECT 5.19 2.42 5.47 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.18 -0.12 1.46 0.83 ;
        RECT 5.285 -0.12 5.475 0.875 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.64 3.19 2.43 ;
        RECT 3 2 3.24 2.43 ;
        RECT 3 0.64 4.02 0.83 ;
        RECT 2.04 2.24 4.02 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.265 0.595 0.455 1.28 ;
      RECT 0.21 1.09 2.695 1.28 ;
      RECT 0.21 1.09 0.4 2.455 ;
      RECT 0.21 2.265 0.55 2.455 ;
      RECT 4.33 0.64 4.61 0.83 ;
      RECT 3.44 1.805 4.52 1.995 ;
      RECT 4.33 0.64 4.52 2.43 ;
      RECT 4.33 2.24 4.61 2.43 ;
  END
END NAND3BBV1_7TV50

MACRO NAND3BBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BBV2_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.26 1.41 8.545 1.92 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.88 1.545 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.03 1.8 1.415 ;
        RECT 1.52 1.225 2.63 1.415 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.04 2.49 1.32 3.48 ;
        RECT 2.715 2.795 3.03 3.48 ;
        RECT 3.635 2.795 3.915 3.48 ;
        RECT 5.335 2.795 5.615 3.48 ;
        RECT 7.04 2.405 7.32 3.48 ;
        RECT 8.635 2.405 8.915 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 -0.12 1.355 0.83 ;
        RECT 2.875 -0.12 3.155 0.635 ;
        RECT 8.685 -0.12 8.965 0.645 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.52 5.64 1.84 ;
        RECT 5.45 1.055 5.64 2.56 ;
        RECT 1.89 2.37 6.47 2.56 ;
        RECT 6.235 0.71 6.515 1.27 ;
        RECT 5.45 1.055 6.515 1.27 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 3.6 -0.24 7.51 1.53 ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.6 3.94 ;
        RECT 7.51 1.46 9.7 3.94 ;
        RECT -0.58 1.53 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.02 0.595 2.21 1.025 ;
      RECT 4.435 0.71 4.715 1.025 ;
      RECT 2.02 0.835 4.715 1.025 ;
      RECT 0.21 1.82 5.195 2.01 ;
      RECT 0.21 0.595 0.4 2.605 ;
      RECT 3.475 0.32 7.43 0.51 ;
      RECT 3.475 0.32 3.755 0.565 ;
      RECT 5.335 0.32 5.615 0.565 ;
      RECT 7.24 0.32 7.43 0.61 ;
      RECT 6.665 1.875 8.02 2.065 ;
      RECT 7.83 0.51 8.02 2.545 ;
  END
END NAND3BBV2_7TV50

MACRO NAND3BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BV1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.96 1.995 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.235 1.56 2.8 1.97 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.46 1.475 1.84 1.855 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 2.445 1.335 3.48 ;
        RECT 2.755 2.79 3.035 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.815 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.605 0.58 3.795 2.48 ;
        RECT 3.44 2.04 3.795 2.48 ;
        RECT 1.905 2.29 3.885 2.48 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.06 3.31 1.25 ;
      RECT 0.2 0.56 0.39 2.48 ;
  END
END NAND3BV1_7TV50

MACRO NAND3BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BV2_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.04 5.91 1.36 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.52 1.8 2.035 ;
        RECT 1.52 1.52 4.4 1.715 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.77 1.08 5.065 1.27 ;
        RECT 4.39 1.08 5.065 1.32 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.795 0.475 3.48 ;
        RECT 1.895 2.795 2.175 3.48 ;
        RECT 3.645 2.795 3.925 3.48 ;
        RECT 5.345 2.795 5.625 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.185 -0.12 0.465 0.49 ;
        RECT 5.295 -0.12 5.575 0.735 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.17 0.69 0.36 2.56 ;
        RECT 0.12 2 0.36 2.56 ;
        RECT 2.84 0.595 3.03 0.88 ;
        RECT 0.17 0.69 3.03 0.88 ;
        RECT 0.12 2.37 4.775 2.56 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 6.275 0.595 6.465 2.11 ;
      RECT 3.255 1.92 6.465 2.11 ;
      RECT 6.24 1.92 6.435 2.52 ;
  END
END NAND3BV2_7TV50

MACRO NAND3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 1.065 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.075 1.76 1.38 ;
        RECT 1.425 1.08 1.905 1.38 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.28 1.04 2.76 1.36 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.765 1.285 3.48 ;
        RECT 2.705 2.385 2.985 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.655 -0.12 2.935 0.595 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2 0.595 0.39 2.43 ;
        RECT 0.12 2 0.39 2.43 ;
        RECT 0.12 2.24 2.135 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
END NAND3V1_7TV50

MACRO NAND3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 0.925 2.89 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.74 1.555 1.035 1.8 ;
        RECT 3.245 1.555 3.555 1.8 ;
        RECT 0.74 1.56 3.555 1.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.695 1.56 5.275 1.84 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.28 2.78 0.56 3.48 ;
        RECT 1.98 2.78 2.26 3.48 ;
        RECT 3.69 2.78 3.97 3.48 ;
        RECT 5.39 2.36 5.67 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.7 -0.12 4.98 0.595 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.33 0.975 0.52 2.55 ;
        RECT 0.12 2 0.52 2.55 ;
        RECT 2.04 0.71 2.32 1.165 ;
        RECT 0.33 0.975 2.32 1.165 ;
        RECT 0.12 2.36 4.82 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.08 -0.24 2.96 1.53 ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.08 3.94 ;
        RECT 2.96 1.46 6.82 3.94 ;
        RECT -0.58 1.53 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.325 0.32 4.035 0.51 ;
      RECT 0.325 0.32 0.515 0.625 ;
      RECT 3.845 0.32 4.035 0.99 ;
      RECT 5.645 0.58 5.835 0.99 ;
      RECT 3.845 0.8 5.835 0.99 ;
  END
END NAND3V2_7TV50

MACRO NAND4BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BV1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 1.055 1.84 ;
        RECT 0.865 1.52 1.055 1.945 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 1.515 3.815 1.945 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.56 2.9 1.915 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.955 1.9 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.295 2.39 1.575 3.48 ;
        RECT 2.995 2.78 3.275 3.48 ;
        RECT 4.695 2.78 4.975 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.345 -0.12 1.625 0.845 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.69 0.595 4.88 2.545 ;
        RECT 4.69 2 5.16 2.545 ;
        RECT 2.145 2.355 5.16 2.545 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.49 0.595 0.68 1.28 ;
      RECT 0.21 1.09 4.4 1.28 ;
      RECT 0.21 1.09 0.4 2.435 ;
      RECT 0.21 2.245 0.725 2.435 ;
  END
END NAND4BV1_7TV50

MACRO NAND4BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BV2_7TV50 0 0 ;
  SIZE 9.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.14 1.04 8.52 1.44 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.705 1.795 1.895 2.19 ;
        RECT 5.805 1.52 6.12 2.19 ;
        RECT 1.705 2 6.12 2.19 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 1.08 2.67 1.8 ;
        RECT 2.48 1.555 2.8 1.8 ;
        RECT 2.48 1.61 5.24 1.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.26 1.125 4.72 1.315 ;
        RECT 4.28 1.08 4.72 1.36 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.335 2.795 0.615 3.48 ;
        RECT 2.035 2.795 2.315 3.48 ;
        RECT 3.735 2.795 4.015 3.48 ;
        RECT 5.435 2.795 5.715 3.48 ;
        RECT 7.135 2.78 7.415 3.48 ;
        RECT 0 3.24 9.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.695 -0.12 3.975 0.49 ;
        RECT 8.615 -0.12 8.895 0.58 ;
        RECT 0 -0.12 9.12 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.375 0.595 0.57 2.32 ;
        RECT 0.12 2 0.57 2.32 ;
        RECT 0.38 0.595 0.57 2.59 ;
        RECT 6.375 0.71 6.565 2.59 ;
        RECT 0.38 2.4 6.565 2.59 ;
        RECT 6.375 0.71 7.395 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 6.75 -0.24 8.195 1.53 ;
        RECT -0.12 -0.24 9.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.75 3.94 ;
        RECT 8.195 1.46 9.7 3.94 ;
        RECT -0.58 1.53 9.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 4.4 0.32 7.94 0.51 ;
      RECT 4.4 0.32 4.59 0.88 ;
      RECT 0.855 0.69 4.59 0.88 ;
      RECT 0.855 0.69 1.045 1.31 ;
      RECT 6.765 1.145 7.94 1.335 ;
      RECT 7.75 0.32 7.94 2.5 ;
      RECT 7.75 2.31 8.265 2.5 ;
  END
END NAND4BV2_7TV50

MACRO NAND4V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.04 3.465 1.415 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.37 1.52 2.76 1.97 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.455 1.03 1.885 1.435 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.52 0.955 1.9 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 2.405 0.575 3.48 ;
        RECT 1.995 2.78 2.275 3.48 ;
        RECT 3.695 2.78 3.975 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.345 -0.12 0.625 0.595 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.69 0.595 3.88 2.55 ;
        RECT 3.69 2 4.2 2.55 ;
        RECT 1.145 2.36 4.2 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
END NAND4V1_7TV50

MACRO NAND4V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.63 1.08 3.28 1.35 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.75 1.555 1.03 1.8 ;
        RECT 0.75 1.56 1.36 1.8 ;
        RECT 3.285 1.555 3.575 1.75 ;
        RECT 0.75 1.56 3.575 1.75 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.315 1.56 4.72 1.81 ;
        RECT 6.78 1.6 7.06 1.81 ;
        RECT 4.315 1.62 7.1 1.81 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.13 1.18 7.16 1.37 ;
        RECT 7.03 1.08 7.6 1.32 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.285 2.78 0.565 3.48 ;
        RECT 1.985 2.78 2.265 3.48 ;
        RECT 3.755 2.78 4.035 3.48 ;
        RECT 5.555 2.78 5.835 3.48 ;
        RECT 7.255 2.405 7.535 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 5.505 -0.12 5.785 0.58 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.17 0.88 0.36 2.55 ;
        RECT 0.12 2 0.36 2.55 ;
        RECT 0.17 0.88 2.235 1.07 ;
        RECT 2.045 0.71 2.325 0.9 ;
        RECT 0.12 2.36 6.685 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.08 -0.24 3.07 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.08 3.94 ;
        RECT 3.07 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.33 0.32 4.04 0.51 ;
      RECT 0.33 0.32 0.52 0.625 ;
      RECT 3.85 0.32 4.04 0.98 ;
      RECT 6.415 0.64 7.485 0.83 ;
      RECT 3.85 0.79 6.605 0.98 ;
  END
END NAND4V2_7TV50

MACRO NAND4XXBBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4XXBBV1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.04 1.99 1.375 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 1.04 0.97 1.41 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.29 1.08 4.72 1.415 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.335 1.56 3.76 1.9 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.13 2.37 2.41 3.48 ;
        RECT 3.88 2.785 4.16 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.38 -0.12 0.66 0.835 ;
        RECT 2.18 -0.12 2.46 0.84 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.68 0.64 5.16 0.83 ;
        RECT 4.92 2 5.16 2.43 ;
        RECT 4.97 0.64 5.16 2.43 ;
        RECT 3.03 2.24 5.16 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.17 0.64 1.56 0.83 ;
      RECT 1.17 0.64 1.36 1.995 ;
      RECT 0.565 1.805 2.785 1.995 ;
      RECT 0.565 1.805 0.76 2.48 ;
  END
END NAND4XXBBV1_7TV50

MACRO NAND4XXBBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4XXBBV2_7TV50 0 0 ;
  SIZE 8.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.48 1.8 1.76 2.32 ;
        RECT 1.48 1.815 1.8 2.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 1.04 0.84 1.36 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.63 1.56 6.16 2.065 ;
        RECT 5.63 1.875 6.76 2.065 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.39 1.17 4.72 1.8 ;
        RECT 4.39 1.17 7.48 1.36 ;
        RECT 7.2 1.17 7.48 1.51 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.855 2.685 2.135 3.48 ;
        RECT 3.555 2.74 3.835 3.48 ;
        RECT 5.24 2.735 5.57 3.48 ;
        RECT 6.94 2.735 7.27 3.48 ;
        RECT 0 3.24 8.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.585 ;
        RECT 1.955 -0.12 2.235 0.585 ;
        RECT 3.755 -0.12 4.035 0.565 ;
        RECT 0 -0.12 8.64 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.105 0.71 7.87 0.9 ;
        RECT 7.32 2 7.87 2.535 ;
        RECT 7.68 0.71 7.87 2.535 ;
        RECT 2.705 2.345 7.87 2.535 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 5.8 -0.24 6.695 1.53 ;
        RECT -0.12 -0.24 8.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.8 3.94 ;
        RECT 6.695 1.46 9.22 3.94 ;
        RECT -0.58 1.53 9.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.08 0.415 1.29 1.345 ;
      RECT 1.08 1.155 3.51 1.345 ;
      RECT 1.08 0.415 1.27 1.895 ;
      RECT 0.3 1.705 1.27 1.895 ;
      RECT 0.3 1.705 0.49 2.475 ;
      RECT 4.39 0.32 8.24 0.51 ;
      RECT 8.05 0.32 8.24 0.61 ;
      RECT 2.9 0.58 3.09 0.955 ;
      RECT 4.39 0.32 4.58 0.955 ;
      RECT 2.9 0.765 4.58 0.955 ;
  END
END NAND4XXBBV2_7TV50

MACRO NOR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2V1_7TV50 0 0 ;
  SIZE 2.4 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.415 1.52 1.8 1.905 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.535 1.03 0.865 1.47 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.355 0.485 3.48 ;
        RECT 0 3.24 2.4 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.61 ;
        RECT 1.955 -0.12 2.235 0.565 ;
        RECT 0 -0.12 2.4 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.595 1.29 0.955 ;
        RECT 1.1 0.765 2.23 0.955 ;
        RECT 2.04 0.765 2.23 2.475 ;
        RECT 2.01 2.195 2.23 2.475 ;
        RECT 2.04 1.52 2.28 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.52 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.98 3.94 ;
    END
  END VNW
END NOR2V1_7TV50

MACRO NOR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.045 1.98 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.84 1.56 1.36 1.8 ;
        RECT 3.2 1.47 3.39 1.75 ;
        RECT 0.84 1.56 3.39 1.75 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.53 2.345 0.81 3.48 ;
        RECT 3.73 2.75 4.01 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.16 -0.12 0.44 0.61 ;
        RECT 2.02 -0.12 2.3 0.39 ;
        RECT 3.88 -0.12 4.16 0.61 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.06 0.61 3.26 0.8 ;
        RECT 3.07 0.61 3.26 1.17 ;
        RECT 3.07 0.98 3.88 1.17 ;
        RECT 3.44 2 3.88 2.43 ;
        RECT 3.69 0.98 3.88 2.43 ;
        RECT 2.13 2.24 3.88 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
END NOR2V2_7TV50

MACRO NOR2V3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2V3_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4 1.17 4.56 1.36 ;
        RECT 4.37 1.17 4.56 1.8 ;
        RECT 4.37 1.56 4.72 1.8 ;
        RECT 4.37 1.61 5.135 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.3 1.8 ;
        RECT 0.75 1.61 3.58 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.275 2.36 0.555 3.48 ;
        RECT 3.73 2.795 4.01 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.27 -0.12 0.46 0.61 ;
        RECT 2.025 -0.12 2.305 0.565 ;
        RECT 3.825 -0.12 4.105 0.565 ;
        RECT 5.625 -0.12 5.905 0.565 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.17 0.595 1.36 0.955 ;
        RECT 2.97 0.595 3.16 0.955 ;
        RECT 4.77 0.595 5.25 0.955 ;
        RECT 1.17 0.765 5.575 0.955 ;
        RECT 5.37 0.765 5.575 2.48 ;
        RECT 2.025 2.29 5.575 2.48 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
END NOR2V3_7TV50

MACRO NOR2V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2V4_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.275 1.84 1.8 ;
        RECT 1.52 1.275 5.41 1.465 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.825 1.695 1.015 2.28 ;
        RECT 0.825 2 1.36 2.28 ;
        RECT 2.22 1.795 2.41 2.19 ;
        RECT 0.825 2 2.41 2.19 ;
        RECT 2.22 1.795 7.095 1.985 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.405 2.36 0.64 3.48 ;
        RECT 3.765 2.795 4.045 3.48 ;
        RECT 7.35 2.735 7.63 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 -0.12 0.535 0.625 ;
        RECT 2.055 -0.12 2.335 0.58 ;
        RECT 3.855 -0.12 4.135 0.58 ;
        RECT 5.715 -0.12 5.995 0.58 ;
        RECT 7.58 -0.12 7.86 0.58 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.2 0.595 1.39 0.975 ;
        RECT 2.105 2.52 2.985 2.71 ;
        RECT 2.48 2.52 2.985 2.76 ;
        RECT 3 0.595 3.19 0.975 ;
        RECT 4.8 0.585 4.99 0.975 ;
        RECT 6.72 0.585 6.91 0.975 ;
        RECT 1.2 0.785 7.495 0.975 ;
        RECT 2.79 2.345 7.495 2.535 ;
        RECT 7.305 0.785 7.495 2.535 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
END NOR2V4_7TV50

MACRO NOR2XBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2XBV1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.8 1.465 1.32 1.655 ;
        RECT 1.08 1.465 1.32 1.88 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.35 1.485 2.76 1.84 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 2.39 1.335 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.83 ;
        RECT 2.855 -0.12 3.135 0.58 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 0.595 2.19 1.21 ;
        RECT 2 1.02 3.19 1.21 ;
        RECT 3 1.02 3.19 2.43 ;
        RECT 3 2 3.24 2.43 ;
        RECT 2.655 2.24 3.24 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.075 1.715 1.265 ;
      RECT 0.2 0.595 0.39 2.43 ;
      RECT 0.2 2.24 0.5 2.43 ;
  END
END NOR2XBV1_7TV50

MACRO NOR2XBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2XBV2_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.84 1.08 1.36 1.37 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.47 1.37 2.775 1.845 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.205 2.68 1.485 3.48 ;
        RECT 4.45 2.745 4.73 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.205 -0.12 1.485 0.635 ;
        RECT 3.005 -0.12 3.285 0.58 ;
        RECT 4.805 -0.12 5.085 0.585 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.15 0.595 2.34 0.97 ;
        RECT 3 0.78 3.24 1.365 ;
        RECT 3.05 0.78 3.24 2.43 ;
        RECT 2.8 2.24 3.24 2.43 ;
        RECT 3.95 0.595 4.14 0.97 ;
        RECT 2.15 0.78 4.14 0.97 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.35 1.805 2.22 1.995 ;
      RECT 3.665 1.805 4.21 1.995 ;
      RECT 0.35 0.595 0.54 2.47 ;
      RECT 0.35 2.28 0.635 2.47 ;
      RECT 2.03 1.805 2.22 2.88 ;
      RECT 3.665 1.805 3.855 2.88 ;
      RECT 2.03 2.69 3.855 2.88 ;
  END
END NOR2XBV2_7TV50

MACRO NOR3BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BV1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 1.52 3.72 1.995 ;
        RECT 3.12 1.805 3.72 1.995 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.46 1.485 1.8 1.995 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.485 1.52 2.76 1.995 ;
        RECT 2.21 1.805 2.76 1.995 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.585 2.78 2.865 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.135 -0.12 1.415 0.565 ;
        RECT 2.935 -0.12 3.215 0.82 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.28 0.58 0.47 2.475 ;
        RECT 0.28 0.795 0.84 1.36 ;
        RECT 2.08 0.58 2.27 0.985 ;
        RECT 0.28 0.795 2.27 0.985 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.835 0.625 4.115 0.815 ;
      RECT 0.755 1.76 0.945 2.43 ;
      RECT 3.925 0.625 4.115 2.43 ;
      RECT 0.755 2.24 4.115 2.43 ;
  END
END NOR3BV1_7TV50

MACRO NOR3BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BV2_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.52 5.64 2.06 ;
        RECT 5.4 1.87 5.895 2.06 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.465 1.51 1.86 1.805 ;
        RECT 1.465 1.615 4.33 1.805 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.795 1.785 0.985 2.28 ;
        RECT 0.795 2.04 1.41 2.28 ;
        RECT 4.81 1.785 5 2.28 ;
        RECT 0.795 2.09 5 2.28 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 2.87 0.495 3.48 ;
        RECT 5.14 2.78 5.42 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.635 ;
        RECT 1.955 -0.12 2.235 0.635 ;
        RECT 3.815 -0.12 4.095 0.44 ;
        RECT 5.675 -0.12 5.96 0.75 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.405 0.96 0.595 2.67 ;
        RECT 1.08 0.54 1.32 1.15 ;
        RECT 2.715 0.64 2.905 1.15 ;
        RECT 0.405 0.96 2.905 1.15 ;
        RECT 0.405 2.48 3.015 2.67 ;
        RECT 2.715 0.64 5.055 0.83 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 6.62 0.595 6.81 1.32 ;
      RECT 3.38 1.13 6.81 1.32 ;
      RECT 3.38 1.13 3.66 1.415 ;
      RECT 6.095 1.13 6.285 2.575 ;
      RECT 5.99 2.385 6.285 2.575 ;
  END
END NOR3BV2_7TV50

MACRO NOR3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.45 1.56 2.71 2.04 ;
        RECT 2.45 1.56 2.8 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.49 1.52 1.835 1.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.84 1.995 ;
        RECT 0.6 1.805 1.085 1.995 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.43 2.4 0.71 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 -0.12 1.405 0.58 ;
        RECT 2.925 -0.12 3.205 0.58 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.27 0.595 0.46 1.045 ;
        RECT 2.07 0.595 2.26 1.045 ;
        RECT 0.27 0.855 3.24 1.045 ;
        RECT 3 0.855 3.24 1.37 ;
        RECT 3.05 0.855 3.24 2.43 ;
        RECT 2.78 2.24 3.24 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
END NOR3V1_7TV50

MACRO NOR3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.485 3.76 1.8 ;
        RECT 3.23 1.485 4.16 1.675 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.375 1.76 2.565 2.2 ;
        RECT 4.4 2.01 4.72 2.28 ;
        RECT 4.875 1.76 5.065 2.2 ;
        RECT 2.375 2.01 5.065 2.2 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.56 1.36 1.995 ;
        RECT 0.63 1.805 1.66 1.995 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.79 1.285 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.585 ;
        RECT 1.955 -0.12 2.235 0.58 ;
        RECT 3.755 -0.12 4.035 0.58 ;
        RECT 5.555 -0.12 5.835 0.585 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.1 0.595 1.29 0.97 ;
        RECT 1.93 0.78 2.12 2.59 ;
        RECT 1.93 0.78 2.28 1.365 ;
        RECT 2.9 0.595 3.09 0.97 ;
        RECT 1.93 2.4 3.735 2.59 ;
        RECT 4.7 0.595 4.89 0.97 ;
        RECT 1.1 0.78 4.89 0.97 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.155 2.24 1.71 2.43 ;
      RECT 1.52 2.24 1.71 2.98 ;
      RECT 1.52 2.79 5.335 2.98 ;
  END
END NOR3V2_7TV50

MACRO NOR4V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 1.52 3.72 1.995 ;
        RECT 3.095 1.805 3.72 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.475 1.37 2.76 1.995 ;
        RECT 2.245 1.805 2.76 1.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.495 1.52 1.81 1.995 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.47 0.885 1.995 ;
        RECT 0.6 1.805 1.025 1.995 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.27 2.37 0.55 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.22 -0.12 0.5 0.59 ;
        RECT 2.02 -0.12 2.3 0.58 ;
        RECT 3.82 -0.12 4.1 0.58 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.165 0.595 1.355 1.025 ;
        RECT 2.965 0.595 3.155 1.025 ;
        RECT 1.165 0.835 4.2 1.025 ;
        RECT 3.96 0.835 4.2 1.365 ;
        RECT 4.01 0.835 4.2 2.47 ;
        RECT 3.37 2.28 4.2 2.47 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
END NOR4V1_7TV50

MACRO NOR4V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.36 1.56 5.68 1.995 ;
        RECT 5.04 1.805 5.97 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.52 1.07 7.62 1.26 ;
        RECT 7.27 1.07 7.62 1.32 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.685 1.07 3.76 1.26 ;
        RECT 3.44 1.07 3.76 1.32 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.8 1.995 ;
        RECT 1.56 1.805 2.77 1.995 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.115 2.76 2.395 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.57 ;
        RECT 2.015 -0.12 2.295 0.435 ;
        RECT 3.93 -0.12 4.215 0.435 ;
        RECT 2.015 -0.12 6.135 0.165 ;
        RECT 5.855 -0.12 6.135 0.435 ;
        RECT 7.715 -0.12 8 0.57 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 0.635 4.15 2.43 ;
        RECT 3.96 2 4.68 2.43 ;
        RECT 3.96 2.24 5.595 2.43 ;
        RECT 1.055 0.635 7.095 0.825 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.515 2.24 3.335 2.43 ;
      RECT 3.145 2.24 3.335 2.98 ;
      RECT 3.145 2.79 7.195 2.98 ;
  END
END NOR4V2_7TV50

MACRO NOR4XXBBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4XXBBV1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 0.95 1.93 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.96 1.9 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.52 3.24 2 ;
        RECT 3 1.81 3.43 2 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 1.505 4.28 2 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.265 2.39 0.545 3.48 ;
        RECT 2.025 2.78 2.305 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.965 -0.12 2.245 0.845 ;
        RECT 3.765 -0.12 4.045 0.595 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.91 0.56 3.1 1.035 ;
        RECT 2.91 0.835 4.9 1.035 ;
        RECT 4.44 0.835 4.9 1.36 ;
        RECT 4.71 0.595 4.9 2.435 ;
        RECT 4.375 2.245 4.9 2.435 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.265 0.64 1.35 0.83 ;
      RECT 1.16 1.08 2.62 1.27 ;
      RECT 1.16 0.64 1.35 2.48 ;
  END
END NOR4XXBBV1_7TV50

MACRO NOR4XXBBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4XXBBV2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 1.04 0.875 1.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.82 1.84 2.28 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.83 1.365 5.02 2.04 ;
        RECT 4.83 1.365 5.16 1.84 ;
        RECT 4.83 1.365 7.31 1.555 ;
        RECT 7.03 1.365 7.31 1.585 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.4 1.805 5.64 2.405 ;
        RECT 5.4 1.805 5.87 1.995 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.22 2.4 0.5 3.48 ;
        RECT 1.92 2.78 2.2 3.48 ;
        RECT 3.72 2.78 4 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.92 -0.12 2.2 0.845 ;
        RECT 3.72 -0.12 4 0.635 ;
        RECT 5.86 -0.12 6.14 0.635 ;
        RECT 7.72 -0.12 8 0.635 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.865 0.595 3.055 1.055 ;
        RECT 4.93 0.595 5.12 1.055 ;
        RECT 6.865 0.55 7.055 1.055 ;
        RECT 2.865 0.865 8.04 1.055 ;
        RECT 7.8 0.865 7.99 2.43 ;
        RECT 6.05 2.24 7.99 2.43 ;
        RECT 7.8 0.865 8.04 1.36 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.17 0.64 1.3 0.83 ;
      RECT 1.11 0.64 1.3 2.595 ;
      RECT 1.11 1.075 2.635 1.265 ;
      RECT 1.11 1.075 1.31 2.595 ;
      RECT 2.87 2.245 4.73 2.435 ;
      RECT 4.54 2.245 4.73 2.98 ;
      RECT 4.54 2.79 7.985 2.98 ;
  END
END NOR4XXBBV2_7TV50

MACRO OA112V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA112V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.815 0.92 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.445 1.895 1.875 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.445 1.07 2.88 1.435 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.32 1.47 3.76 1.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.135 2.495 2.415 3.48 ;
        RECT 3.885 2.495 4.165 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.885 -0.12 4.165 0.58 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.83 0.58 5.02 2.595 ;
        RECT 4.83 2 5.16 2.595 ;
        RECT 4.735 2.405 5.16 2.595 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.585 -0.24 2.325 1.555 ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.585 3.94 ;
        RECT 2.325 1.46 5.86 3.94 ;
        RECT -0.58 1.555 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.31 0.32 2.42 0.51 ;
      RECT 0.31 0.32 0.5 0.61 ;
      RECT 2.23 0.32 2.42 0.61 ;
      RECT 1.17 0.71 1.505 0.9 ;
      RECT 1.17 0.71 1.36 2.29 ;
      RECT 4.305 1.75 4.495 2.29 ;
      RECT 0.58 2.1 4.495 2.29 ;
      RECT 0.58 2.1 0.77 2.57 ;
      RECT 3.08 2.1 3.27 2.57 ;
  END
END OA112V1_7TV50

MACRO OA112V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA112V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.975 0.94 1.38 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.8 2.09 ;
        RECT 1.56 1.9 1.94 2.09 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.44 0.98 2.84 1.36 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.56 3.76 2.105 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.135 2.795 2.415 3.48 ;
        RECT 3.885 2.795 4.165 3.48 ;
        RECT 5.685 2.39 5.965 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.885 -0.12 4.165 0.58 ;
        RECT 5.685 -0.12 5.965 0.58 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.83 0.51 5.02 2.64 ;
        RECT 4.83 2 5.16 2.325 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.585 -0.24 2.325 1.555 ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.585 3.94 ;
        RECT 2.325 1.46 6.82 3.94 ;
        RECT -0.58 1.555 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.31 0.32 2.42 0.51 ;
      RECT 0.31 0.32 0.5 0.65 ;
      RECT 2.23 0.32 2.42 0.65 ;
      RECT 1.17 0.71 1.505 0.9 ;
      RECT 1.17 0.71 1.36 2.525 ;
      RECT 4.305 1.75 4.495 2.525 ;
      RECT 0.535 2.335 4.495 2.525 ;
  END
END OA112V2_7TV50

MACRO OA12V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA12V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.8 2.12 ;
        RECT 1.435 1.93 1.8 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 0.84 2.12 ;
        RECT 0.6 1.93 1.05 2.12 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.415 1.56 2.605 2.165 ;
        RECT 2.415 1.56 2.8 1.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 2.48 0.575 3.48 ;
        RECT 2.99 2.475 3.27 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.98 -0.12 3.26 0.875 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.87 0.64 4.2 0.83 ;
        RECT 3.96 2 4.2 2.435 ;
        RECT 4.01 0.64 4.2 2.435 ;
        RECT 3.84 2.245 4.2 2.435 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.665 -0.24 2.655 1.585 ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.665 3.94 ;
        RECT 2.655 1.46 4.9 3.94 ;
        RECT -0.58 1.585 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.565 0.72 2.3 0.91 ;
      RECT 0.205 0.595 0.395 1.265 ;
      RECT 1.565 0.72 1.755 1.265 ;
      RECT 0.205 1.075 1.755 1.265 ;
      RECT 1.105 0.32 2.69 0.51 ;
      RECT 1.105 0.32 1.295 0.875 ;
      RECT 2.5 0.32 2.69 1.3 ;
      RECT 2 1.11 3.67 1.3 ;
      RECT 2 1.11 2.19 2.585 ;
      RECT 1.895 2.395 2.19 2.585 ;
  END
END OA12V1_7TV50

MACRO OA12V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA12V2_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.52 1.8 2.09 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 0.92 1.9 ;
        RECT 0.715 1.56 0.92 2.135 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.415 1.52 2.605 2.135 ;
        RECT 2.415 1.52 2.76 1.84 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.295 2.4 0.575 3.48 ;
        RECT 2.855 2.405 3.135 3.48 ;
        RECT 4.555 2.4 4.835 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.98 -0.12 3.26 0.67 ;
        RECT 4.78 -0.12 5.06 0.57 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.87 0.625 4.2 0.815 ;
        RECT 3.96 2 4.2 2.555 ;
        RECT 4.01 0.625 4.2 2.555 ;
        RECT 3.705 2.365 4.2 2.555 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.385 -0.24 2.605 1.54 ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.385 3.94 ;
        RECT 2.605 1.46 5.86 3.94 ;
        RECT -0.58 1.54 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.565 0.71 2.3 0.9 ;
      RECT 0.205 0.58 0.395 1.265 ;
      RECT 1.565 0.71 1.755 1.265 ;
      RECT 0.205 1.075 1.755 1.265 ;
      RECT 1.105 0.32 2.69 0.51 ;
      RECT 1.105 0.32 1.295 0.86 ;
      RECT 2.5 0.32 2.69 1.32 ;
      RECT 3.355 1.075 3.635 1.32 ;
      RECT 2 1.13 3.635 1.32 ;
      RECT 2 1.13 2.19 2.555 ;
      RECT 1.895 2.365 2.19 2.555 ;
  END
END OA12V2_7TV50

MACRO OA21BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21BV1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.53 1.075 0.9 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.86 2.045 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.52 3.24 1.995 ;
        RECT 3 1.805 3.455 1.995 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.95 2.79 2.23 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.835 ;
        RECT 1.955 -0.12 2.235 0.83 ;
        RECT 3.755 -0.12 4.035 0.58 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9 0.595 3.09 0.97 ;
        RECT 2.9 0.78 3.845 0.97 ;
        RECT 3.48 0.78 3.845 1.36 ;
        RECT 3.655 0.78 3.845 2.43 ;
        RECT 3.55 2.24 3.845 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.1 0.595 1.29 2.435 ;
      RECT 2.47 1.76 2.66 2.435 ;
      RECT 0.29 2.245 2.66 2.435 ;
  END
END OA21BV1_7TV50

MACRO OA21BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21BV2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.4 0.875 1.94 ;
        RECT 0.6 1.66 0.92 1.94 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.87 2.035 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.22 1.56 3.76 1.895 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.995 2.775 2.275 3.48 ;
        RECT 5.21 2.39 5.49 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.25 -0.12 0.53 0.845 ;
        RECT 2.05 -0.12 2.33 0.845 ;
        RECT 3.855 -0.12 4.135 0.58 ;
        RECT 5.655 -0.12 5.935 0.595 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.595 3.19 1.195 ;
        RECT 3.96 1.005 4.2 1.36 ;
        RECT 4.01 1.005 4.2 2.43 ;
        RECT 3.595 2.24 4.2 2.43 ;
        RECT 4.8 0.595 4.99 1.195 ;
        RECT 3 1.005 4.99 1.195 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.17 0.595 1.395 1.32 ;
      RECT 2.425 1.075 2.705 1.32 ;
      RECT 1.17 1.13 2.705 1.32 ;
      RECT 4.445 1.805 5.1 1.995 ;
      RECT 1.17 0.595 1.36 2.43 ;
      RECT 0.31 2.24 2.91 2.43 ;
      RECT 2.72 2.24 2.91 2.82 ;
      RECT 4.445 1.805 4.635 2.82 ;
      RECT 2.72 2.63 4.635 2.82 ;
  END
END OA21BV2_7TV50

MACRO OA221V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.52 3.24 2.12 ;
        RECT 3 1.93 3.435 2.12 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.9 1.52 4.2 2.075 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.56 2.32 2.12 ;
        RECT 2 1.93 2.685 2.12 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.44 0.895 1.8 1.36 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.51 0.84 2.12 ;
        RECT 0.6 1.93 1.01 2.12 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.12 2.755 1.4 3.48 ;
        RECT 4.44 2.755 4.72 3.48 ;
        RECT 5.03 2.795 5.31 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.575 -0.12 3.855 0.815 ;
        RECT 5.375 -0.12 5.655 0.835 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.88 2 6.12 2.435 ;
        RECT 6.32 0.58 6.51 2.435 ;
        RECT 5.88 2.245 6.51 2.435 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.055 -0.24 3.18 1.585 ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.055 3.94 ;
        RECT 3.18 1.46 7.3 3.94 ;
        RECT -0.58 1.585 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.065 0.375 3.275 0.565 ;
      RECT 2.025 0.765 2.405 0.955 ;
      RECT 2.215 0.765 2.405 1.205 ;
      RECT 4.52 0.58 4.71 1.205 ;
      RECT 2.215 1.015 4.71 1.205 ;
      RECT 4.53 1.765 5.64 2.045 ;
      RECT 0.21 0.33 0.4 2.555 ;
      RECT 4.53 1.765 4.72 2.555 ;
      RECT 0.21 2.365 4.72 2.555 ;
  END
END OA221V1_7TV50

MACRO OA221V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221V2_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.52 3.24 2.09 ;
        RECT 3 1.9 3.42 2.09 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.885 1.52 4.2 2.09 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.52 2.34 2.09 ;
        RECT 2.04 1.9 2.465 2.09 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4 0.98 1.8 1.36 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.98 1.01 1.36 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.06 2.795 1.34 3.48 ;
        RECT 4.26 2.755 4.54 3.48 ;
        RECT 5.435 2.4 5.715 3.48 ;
        RECT 7.135 2.38 7.415 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.585 -0.12 3.865 0.66 ;
        RECT 5.385 -0.12 5.665 0.675 ;
        RECT 7.185 -0.12 7.465 0.58 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.33 0.58 6.52 2.48 ;
        RECT 6.33 1.52 6.6 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.03 -0.24 3.155 1.53 ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.03 3.94 ;
        RECT 3.155 1.46 8.26 3.94 ;
        RECT -0.58 1.53 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.12 0.32 3.23 0.51 ;
      RECT 1.12 0.32 1.31 0.61 ;
      RECT 3.04 0.32 3.23 0.61 ;
      RECT 4.14 0.625 4.765 0.815 ;
      RECT 2.035 0.71 2.405 0.9 ;
      RECT 2.215 0.71 2.405 1.205 ;
      RECT 4.14 0.625 4.33 1.205 ;
      RECT 2.215 1.015 4.33 1.205 ;
      RECT 5.805 1.03 5.995 1.835 ;
      RECT 4.79 1.645 5.995 1.835 ;
      RECT 0.21 0.5 0.4 2.53 ;
      RECT 4.79 1.645 4.98 2.53 ;
      RECT 0.21 2.34 4.98 2.53 ;
  END
END OA221V2_7TV50

MACRO OA222V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222V1_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.51 1.03 0.93 1.375 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.455 1.89 1.88 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.43 1.465 2.815 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.32 1.47 3.76 1.8 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.88 1.03 6.18 1.52 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.92 1.465 5.33 1.945 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.38 2.455 0.66 3.48 ;
        RECT 3.715 2.47 3.995 3.48 ;
        RECT 6.32 2.405 6.6 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.485 -0.12 4.765 0.83 ;
        RECT 6.31 -0.12 6.59 0.83 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.21 0.64 7.51 0.83 ;
        RECT 7.32 0.64 7.51 2.435 ;
        RECT 7.17 2.245 7.51 2.435 ;
        RECT 7.32 1.52 7.56 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.58 -0.24 3.605 1.53 ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.58 3.94 ;
        RECT 3.605 1.46 8.26 3.94 ;
        RECT -0.58 1.53 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.17 0.32 4.17 0.51 ;
      RECT 0.17 0.32 0.45 0.83 ;
      RECT 3.89 0.32 4.17 0.83 ;
      RECT 2.075 0.32 2.265 0.875 ;
      RECT 2.93 0.71 3.21 1.235 ;
      RECT 5.43 0.595 5.62 1.235 ;
      RECT 2.93 1.045 5.62 1.235 ;
      RECT 1.13 0.71 1.41 0.9 ;
      RECT 6.74 1.765 6.93 2.065 ;
      RECT 5.93 1.875 6.93 2.065 ;
      RECT 1.13 0.71 1.32 2.285 ;
      RECT 1.13 2.08 4.475 2.27 ;
      RECT 1.13 2.08 2.23 2.285 ;
      RECT 4.285 2.08 4.475 2.56 ;
      RECT 5.93 1.875 6.12 2.56 ;
      RECT 4.285 2.37 6.12 2.56 ;
      RECT 2.04 2.08 2.23 2.61 ;
  END
END OA222V1_7TV50

MACRO OA222V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222V2_7TV50 0 0 ;
  SIZE 8.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.03 0.92 1.5 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.04 1.935 1.44 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.43 1.465 2.815 1.99 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.275 1.56 3.76 1.99 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.31 1.52 5.64 2 ;
        RECT 5.31 1.81 5.765 2 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.34 1.52 4.68 2.005 ;
        RECT 4.34 1.81 4.955 2.005 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.47 2.4 0.75 3.48 ;
        RECT 3.67 2.775 3.95 3.48 ;
        RECT 5.86 2.78 6.14 3.48 ;
        RECT 7.56 2.78 7.84 3.48 ;
        RECT 0 3.24 8.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.485 -0.12 4.765 0.645 ;
        RECT 6.285 -0.12 6.565 0.645 ;
        RECT 8.085 -0.12 8.365 0.595 ;
        RECT 0 -0.12 8.64 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.23 0.595 7.42 2.545 ;
        RECT 6.71 2.355 7.42 2.545 ;
        RECT 7.23 2 7.56 2.32 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.58 -0.24 3.605 1.53 ;
        RECT -0.12 -0.24 8.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.58 3.94 ;
        RECT 3.605 1.46 9.22 3.94 ;
        RECT -0.58 1.53 9.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.215 0.32 4.13 0.51 ;
      RECT 0.215 0.32 0.405 0.75 ;
      RECT 2.03 0.32 2.31 0.83 ;
      RECT 3.94 0.32 4.13 0.845 ;
      RECT 2.91 0.71 3.21 0.9 ;
      RECT 3.02 0.71 3.21 1.235 ;
      RECT 5.43 0.595 5.62 1.235 ;
      RECT 3.02 1.045 5.62 1.235 ;
      RECT 1.13 0.71 1.41 0.9 ;
      RECT 5.965 1.075 6.94 1.265 ;
      RECT 1.13 0.71 1.32 2.5 ;
      RECT 5.965 1.075 6.155 2.5 ;
      RECT 1.13 2.31 6.155 2.5 ;
  END
END OA222V2_7TV50

MACRO OA22V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.425 1.445 2.805 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.405 1.52 3.72 1.98 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.44 1.845 1.8 2.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.48 0.945 1.8 ;
        RECT 0.755 1.48 0.945 2.15 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.335 2.485 0.615 3.48 ;
        RECT 4.195 2.395 4.48 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.565 ;
        RECT 4.47 -0.12 4.75 0.57 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.43 0.58 5.62 2.475 ;
        RECT 5.4 1.04 5.64 1.36 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.345 -0.24 3.755 1.535 ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.345 3.94 ;
        RECT 3.755 1.46 6.82 3.94 ;
        RECT -0.58 1.535 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2 0.32 4.11 0.51 ;
      RECT 3.92 0.32 4.11 0.61 ;
      RECT 0.2 0.33 0.39 0.955 ;
      RECT 2 0.32 2.19 0.955 ;
      RECT 0.2 0.765 2.19 0.955 ;
      RECT 2.915 0.71 3.195 1.25 ;
      RECT 2.915 1.06 5.14 1.25 ;
      RECT 3.005 0.71 3.195 2.675 ;
      RECT 1.935 2.485 3.195 2.675 ;
  END
END OA22V1_7TV50

MACRO OA22V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22V2_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.425 1.445 2.805 1.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.405 1.52 3.735 1.98 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.44 1.52 1.8 1.92 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.425 0.945 1.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.335 2.4 0.615 3.48 ;
        RECT 3.9 2.79 4.24 3.48 ;
        RECT 6.285 2.4 6.565 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.565 ;
        RECT 4.47 -0.12 4.75 0.57 ;
        RECT 6.285 -0.12 6.565 0.565 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.43 0.43 5.62 2.68 ;
        RECT 5.4 1.52 5.64 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.345 -0.24 3.755 1.535 ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.345 3.94 ;
        RECT 3.755 1.46 7.3 3.94 ;
        RECT -0.58 1.535 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2 0.32 4.155 0.51 ;
      RECT 3.845 0.32 4.155 0.565 ;
      RECT 0.2 0.495 0.39 0.955 ;
      RECT 2 0.32 2.19 0.955 ;
      RECT 0.2 0.765 2.19 0.955 ;
      RECT 2.915 0.71 3.195 1.035 ;
      RECT 2.915 0.845 4.895 1.035 ;
      RECT 4.705 0.845 4.895 2.41 ;
      RECT 2.035 2.22 4.895 2.41 ;
      RECT 2.035 2.22 2.315 2.52 ;
  END
END OA22V2_7TV50

MACRO OA31V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.56 1.875 1.99 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.495 1.52 2.8 1.995 ;
        RECT 2.18 1.805 2.8 1.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.38 1.075 3.76 1.465 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.555 1.52 0.84 2.04 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.385 0.485 3.48 ;
        RECT 3.47 2.66 3.75 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.955 -0.12 2.235 0.82 ;
        RECT 3.755 -0.12 4.035 0.83 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 2 4.89 2.43 ;
        RECT 4.7 0.595 4.89 2.43 ;
        RECT 4.32 2.24 4.89 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.055 0.63 1.75 0.82 ;
      RECT 2.68 0.63 3.135 0.82 ;
      RECT 1.56 0.63 1.75 1.225 ;
      RECT 2.68 0.63 2.87 1.225 ;
      RECT 1.56 1.035 2.87 1.225 ;
      RECT 0.2 0.595 0.39 1.32 ;
      RECT 0.2 1.13 1.245 1.32 ;
      RECT 1.055 1.13 1.245 2.43 ;
      RECT 3.925 1.76 4.115 2.43 ;
      RECT 1.055 2.24 4.115 2.43 ;
  END
END OA31V1_7TV50

MACRO OA31V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.425 1.905 2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.31 1.56 2.59 2 ;
        RECT 2.31 1.56 2.8 1.81 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.38 1.075 3.76 1.46 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.5 1.56 0.88 2.045 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.23 2.345 0.515 3.48 ;
        RECT 3.435 2.725 3.715 3.48 ;
        RECT 5.135 2.75 5.415 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.045 -0.12 2.325 0.39 ;
        RECT 3.905 -0.12 4.185 0.625 ;
        RECT 5.705 -0.12 5.985 0.61 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.85 0.595 5.04 1.495 ;
        RECT 4.85 1.305 5.655 1.495 ;
        RECT 5.4 2 5.655 2.535 ;
        RECT 5.465 1.305 5.655 2.535 ;
        RECT 4.285 2.345 5.655 2.535 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.085 0.59 3.285 0.78 ;
      RECT 0.23 0.58 0.42 1.17 ;
      RECT 0.23 0.98 1.32 1.17 ;
      RECT 3.53 1.81 4.94 2 ;
      RECT 1.085 0.98 1.32 2.44 ;
      RECT 3.53 1.81 3.72 2.44 ;
      RECT 1.085 2.25 3.72 2.44 ;
  END
END OA31V2_7TV50

MACRO OA32V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA32V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.5 2.28 1.98 ;
        RECT 2.04 1.755 2.41 1.98 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.52 3.36 1.93 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.865 1.47 4.2 1.925 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.33 2 1.61 2.39 ;
        RECT 1.33 2 1.8 2.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.12 2 0.36 2.39 ;
        RECT 0.12 2.2 0.86 2.39 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.78 0.485 3.48 ;
        RECT 4.155 2.78 4.435 3.48 ;
        RECT 4.745 2.395 5.025 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.83 ;
        RECT 5.365 -0.12 5.6 0.625 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.88 2 6.12 2.44 ;
        RECT 5.93 0.64 6.12 2.44 ;
        RECT 5.595 2.24 6.12 2.44 ;
        RECT 5.93 0.64 6.545 0.83 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.125 -0.24 3.76 1.85 ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.125 3.94 ;
        RECT 3.76 1.46 7.3 3.94 ;
        RECT -0.58 1.85 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.955 0.64 4.155 0.83 ;
      RECT 0.2 0.595 0.39 1.22 ;
      RECT 1.955 0.64 2.145 1.22 ;
      RECT 0.2 1.03 2.145 1.22 ;
      RECT 4.82 0.595 5.01 1.28 ;
      RECT 2.61 1.03 5.01 1.22 ;
      RECT 4.82 1.09 5.72 1.28 ;
      RECT 2.61 1.03 2.8 2.835 ;
      RECT 1.805 2.645 2.8 2.835 ;
  END
END OA32V1_7TV50

MACRO OA32V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA32V2_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.52 2.405 1.84 ;
        RECT 2.215 1.52 2.405 2.05 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.52 3.36 2.005 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 1.52 4.2 2.005 ;
        RECT 3.735 1.765 4.2 2.005 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.52 1.32 2.06 ;
        RECT 1.08 1.87 1.61 2.06 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.12 1.52 0.36 2.06 ;
        RECT 0.12 1.87 0.86 2.06 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.205 2.395 0.485 3.48 ;
        RECT 4.21 2.4 4.49 3.48 ;
        RECT 5.415 2.4 5.695 3.48 ;
        RECT 7.115 2.405 7.395 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.605 ;
        RECT 5.365 -0.12 5.645 0.6 ;
        RECT 7.165 -0.12 7.445 0.59 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.31 0.595 6.5 2.48 ;
        RECT 6.31 2 6.6 2.325 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.125 -0.24 3.705 1.525 ;
        RECT 2.8 -0.24 3.705 1.535 ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.125 3.94 ;
        RECT -0.58 1.525 2.8 3.94 ;
        RECT 3.705 1.46 8.26 3.94 ;
        RECT -0.58 1.535 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2 0.32 4.11 0.51 ;
      RECT 3.92 0.32 4.11 0.65 ;
      RECT 0.2 0.54 0.39 0.995 ;
      RECT 2 0.32 2.19 0.995 ;
      RECT 0.2 0.805 2.19 0.995 ;
      RECT 2.915 0.71 3.195 1.265 ;
      RECT 4.82 0.54 5.01 1.265 ;
      RECT 2.605 1.075 6.02 1.265 ;
      RECT 2.605 1.075 2.795 2.835 ;
      RECT 1.805 2.645 2.795 2.835 ;
  END
END OA32V2_7TV50

MACRO OA33V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33V1_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.405 1.56 2.595 2.11 ;
        RECT 2.405 1.56 2.8 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.845 2.11 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 0.97 1.8 ;
        RECT 0.78 1.56 0.97 2.11 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.25 1.465 3.72 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 1.52 4.2 2.13 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.795 1.52 5.275 1.84 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.385 2.455 0.665 3.48 ;
        RECT 5.145 2.78 5.425 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.875 -0.12 4.155 0.83 ;
        RECT 5.675 -0.12 5.955 0.845 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.36 2 6.81 2.435 ;
        RECT 6.62 0.595 6.81 2.435 ;
        RECT 5.995 2.245 6.81 2.435 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.595 -0.24 3.7 1.53 ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.595 3.94 ;
        RECT 3.7 1.46 7.78 3.94 ;
        RECT -0.58 1.53 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.055 0.32 3.21 0.51 ;
      RECT 1.055 0.32 1.335 0.83 ;
      RECT 3.02 0.32 3.21 1.22 ;
      RECT 4.82 0.595 5.01 1.22 ;
      RECT 3.02 1.03 5.01 1.22 ;
      RECT 2.015 0.71 2.295 0.9 ;
      RECT 0.2 0.595 0.39 1.22 ;
      RECT 2.015 0.71 2.205 1.22 ;
      RECT 0.2 1.03 2.205 1.22 ;
      RECT 5.565 1.445 5.755 2.3 ;
      RECT 4.685 2.11 5.755 2.3 ;
      RECT 1.17 1.03 1.36 2.605 ;
      RECT 4.685 2.11 4.875 2.605 ;
      RECT 1.17 2.415 4.875 2.605 ;
  END
END OA33V1_7TV50

MACRO OA33V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 1.45 2.89 1.84 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.925 1.915 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.46 1.515 0.975 1.815 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.415 1.5 3.805 1.93 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.395 1.505 4.705 1.97 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.265 1.52 5.64 1.905 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.52 2.405 0.8 3.48 ;
        RECT 5.575 2.795 5.855 3.48 ;
        RECT 7.275 2.405 7.555 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.975 -0.12 4.255 0.7 ;
        RECT 5.775 -0.12 6.055 0.7 ;
        RECT 7.575 -0.12 7.855 0.635 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.72 0.595 6.91 2.555 ;
        RECT 6.425 2.365 6.91 2.555 ;
        RECT 6.72 1.56 7.12 1.8 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.21 -0.24 3.075 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.21 3.94 ;
        RECT 3.075 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.155 0.32 3.31 0.51 ;
      RECT 1.155 0.32 1.435 0.7 ;
      RECT 3.12 0.32 3.31 1.09 ;
      RECT 4.92 0.595 5.11 1.09 ;
      RECT 3.12 0.9 5.11 1.09 ;
      RECT 0.3 0.595 0.49 1.09 ;
      RECT 2.115 0.71 2.395 1.09 ;
      RECT 0.3 0.9 2.395 1.09 ;
      RECT 2.125 0.71 2.315 2.555 ;
      RECT 5.995 1.765 6.185 2.555 ;
      RECT 2.125 2.365 6.185 2.555 ;
  END
END OA33V2_7TV50

MACRO OAI211V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.445 1.52 2.895 1.845 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.39 1.52 3.84 1.845 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.015 1.04 1.32 1.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 2.01 1.845 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.265 2.795 1.545 3.48 ;
        RECT 3.715 2.405 3.995 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.965 -0.12 3.245 0.58 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.365 0.64 0.65 0.83 ;
        RECT 0.12 1.52 0.65 1.84 ;
        RECT 0.46 0.64 0.65 2.55 ;
        RECT 0.46 2.36 2.395 2.55 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.11 0.595 2.3 0.97 ;
      RECT 3.91 0.595 4.1 0.97 ;
      RECT 2.11 0.78 4.1 0.97 ;
  END
END OAI211V1_7TV50

MACRO OAI211V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.88 1.52 6.12 2.035 ;
        RECT 5.175 1.845 6.225 2.035 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.435 1.08 4.625 1.36 ;
        RECT 4.88 1.08 5.2 1.32 ;
        RECT 4.435 1.08 7.315 1.27 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.08 1.36 1.32 ;
        RECT 1.04 1.1 2.575 1.29 ;
        RECT 2.385 1.1 2.575 1.38 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 1.56 3.28 1.8 ;
        RECT 0.615 1.61 3.48 1.8 ;
        RECT 3.29 1.61 3.48 2.11 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.615 0.435 3.48 ;
        RECT 1.915 2.7 2.195 3.48 ;
        RECT 3.855 2.795 4.135 3.48 ;
        RECT 7.225 2.405 7.505 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.68 -0.12 4.96 0.39 ;
        RECT 6.6 -0.12 6.88 0.39 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.965 0.71 3.56 0.9 ;
        RECT 3.37 0.71 3.56 1.215 ;
        RECT 3.37 1.025 4.2 1.215 ;
        RECT 3.96 1.52 4.2 1.84 ;
        RECT 4.01 1.025 4.2 2.5 ;
        RECT 1.005 2.31 5.85 2.5 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.195 -0.24 3.6 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.195 3.94 ;
        RECT 3.6 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.25 0.32 3.955 0.51 ;
      RECT 0.25 0.32 0.44 0.625 ;
      RECT 3.765 0.32 3.955 0.825 ;
      RECT 3.765 0.635 7.84 0.825 ;
  END
END OAI211V2_7TV50

MACRO OAI21BV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BV1_7TV50 0 0 ;
  SIZE 4.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.3 1.04 0.84 1.365 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.905 1.52 3.355 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.865 1.52 4.315 1.84 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.77 2.79 2.05 3.48 ;
        RECT 4.22 2.395 4.5 3.48 ;
        RECT 0 3.24 4.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.83 ;
        RECT 3.455 -0.12 3.735 0.58 ;
        RECT 0 -0.12 4.8 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.655 0.64 2.28 0.83 ;
        RECT 2.04 1.52 2.28 1.84 ;
        RECT 2.09 0.64 2.28 2.43 ;
        RECT 2.09 2.24 2.9 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.11 1.075 1.855 1.265 ;
      RECT 1.11 0.595 1.3 2.46 ;
      RECT 0.86 2.27 1.3 2.46 ;
      RECT 2.6 0.595 2.79 0.97 ;
      RECT 4.4 0.595 4.59 0.97 ;
      RECT 2.6 0.78 4.59 0.97 ;
  END
END OAI21BV1_7TV50

MACRO OAI21BV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21BV2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.875 0.84 2.32 ;
        RECT 0.6 1.875 1.155 2.065 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.84 1.075 6.16 1.32 ;
        RECT 5.315 1.075 6.43 1.265 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.88 1.56 5.2 2.065 ;
        RECT 6.68 1.765 6.87 2.065 ;
        RECT 4.33 1.875 6.87 2.065 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.495 2.79 0.775 3.48 ;
        RECT 2.155 2.405 2.435 3.48 ;
        RECT 3.855 2.795 4.135 3.48 ;
        RECT 7.11 2.405 7.39 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.445 -0.12 0.725 0.615 ;
        RECT 4.815 -0.12 5.095 0.435 ;
        RECT 6.735 -0.12 7.015 0.435 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.895 0.71 3.24 0.9 ;
        RECT 3 1.52 3.24 1.84 ;
        RECT 3.05 0.71 3.24 2.595 ;
        RECT 2.97 2.405 5.79 2.595 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.205 -0.24 3.825 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.205 3.94 ;
        RECT 3.825 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.39 1.875 2.765 2.065 ;
      RECT 2.575 1.83 2.765 2.11 ;
      RECT 1.39 0.55 1.58 2.545 ;
      RECT 1.935 0.32 4.09 0.51 ;
      RECT 1.935 0.32 2.225 0.58 ;
      RECT 3.9 0.32 4.09 0.825 ;
      RECT 3.9 0.635 7.975 0.825 ;
  END
END OAI21BV2_7TV50

MACRO OAI21V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.56 1.84 2.045 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 1 2.045 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.365 1.475 2.76 1.95 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.375 2.405 0.655 3.48 ;
        RECT 2.885 2.795 3.165 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 -0.12 1.405 0.565 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.97 0.58 3.16 2.435 ;
        RECT 1.975 2.245 3.16 2.435 ;
        RECT 2.97 1.52 3.24 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.27 0.58 0.46 0.955 ;
      RECT 2.07 0.58 2.26 0.955 ;
      RECT 0.27 0.765 2.26 0.955 ;
  END
END OAI21V1_7TV50

MACRO OAI21V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.56 2.32 1.8 ;
        RECT 1.53 1.56 2.56 1.75 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.725 1.765 0.915 2.19 ;
        RECT 1.04 2 1.38 2.28 ;
        RECT 3.175 1.765 3.365 2.19 ;
        RECT 0.725 2 3.365 2.19 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.24 1.44 5.68 1.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.305 2.405 0.585 3.48 ;
        RECT 3.505 2.795 3.785 3.48 ;
        RECT 5.205 2.405 5.485 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.565 ;
        RECT 2.855 -0.12 3.135 0.565 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.4 1.56 4.72 1.8 ;
        RECT 4.53 0.71 4.72 2.595 ;
        RECT 1.905 2.405 4.72 2.595 ;
        RECT 4.53 0.71 4.995 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.41 -0.24 5.3 1.545 ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.41 3.94 ;
        RECT 5.3 1.46 6.82 3.94 ;
        RECT -0.58 1.545 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.8 0.32 5.91 0.51 ;
      RECT 5.72 0.32 5.91 0.61 ;
      RECT 0.2 0.58 0.39 0.955 ;
      RECT 2 0.58 2.19 0.955 ;
      RECT 3.8 0.32 3.99 0.955 ;
      RECT 0.2 0.765 3.99 0.955 ;
  END
END OAI21V2_7TV50

MACRO OAI221V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.835 1.52 2.28 1.89 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.975 1.455 1.395 1.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.495 1.505 2.925 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.45 1.52 3.94 1.855 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.92 1.52 5.185 2.07 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.6 2.405 0.88 3.48 ;
        RECT 4.035 2.795 4.315 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.365 -0.12 1.645 0.565 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.75 0.595 5.94 2.555 ;
        RECT 2.3 2.36 5.94 2.555 ;
        RECT 5.75 1.515 6.12 1.845 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.835 -0.24 5.115 1.53 ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.835 3.94 ;
        RECT 5.115 1.46 6.82 3.94 ;
        RECT -0.58 1.53 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.31 0.32 4.465 0.51 ;
      RECT 4.185 0.32 4.465 0.565 ;
      RECT 0.51 0.505 0.7 0.955 ;
      RECT 2.31 0.32 2.5 0.955 ;
      RECT 0.51 0.765 2.5 0.955 ;
      RECT 3.225 0.71 3.505 0.955 ;
      RECT 4.82 0.595 5.01 0.955 ;
      RECT 3.225 0.765 5.01 0.955 ;
  END
END OAI221V1_7TV50

MACRO OAI221V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221V2_7TV50 0 0 ;
  SIZE 10.56 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.96 2.025 2.32 2.28 ;
        RECT 1.96 2.025 2.995 2.215 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.025 1.56 1.36 1.8 ;
        RECT 1.025 1.61 3.8 1.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.265 1.3 8.04 1.49 ;
        RECT 7.68 1.3 8.04 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.37 1.505 4.68 2.08 ;
        RECT 4.37 1.89 7.235 2.08 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.68 1.56 10.32 1.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.685 2.405 0.965 3.48 ;
        RECT 3.995 2.795 4.275 3.48 ;
        RECT 7.505 2.795 7.785 3.48 ;
        RECT 9.365 2.795 9.645 3.48 ;
        RECT 0 3.24 10.56 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.2 -0.12 1.48 0.565 ;
        RECT 3 -0.12 3.28 0.565 ;
        RECT 0 -0.12 10.56 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.34 2.48 3.36 2.67 ;
        RECT 3.205 2.405 9.355 2.595 ;
        RECT 9.135 0.71 9.355 2.595 ;
        RECT 9.135 0.71 9.42 1.37 ;
        RECT 9.135 1.04 9.48 1.37 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 5.335 -0.24 9.78 1.545 ;
        RECT -0.12 -0.24 10.68 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.335 3.94 ;
        RECT 9.78 1.46 11.14 3.94 ;
        RECT -0.58 1.545 11.14 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.345 0.58 0.535 0.955 ;
      RECT 2.145 0.58 2.335 0.955 ;
      RECT 3.945 0.58 4.135 0.995 ;
      RECT 5.76 0.715 6.04 0.995 ;
      RECT 0.345 0.765 4.135 0.955 ;
      RECT 7.56 0.715 7.84 0.995 ;
      RECT 3.945 0.805 7.84 0.995 ;
      RECT 4.8 0.32 10.375 0.51 ;
      RECT 4.8 0.32 5.08 0.565 ;
      RECT 6.66 0.32 6.94 0.565 ;
      RECT 8.175 0.32 8.455 0.565 ;
      RECT 10.095 0.32 10.375 0.565 ;
  END
END OAI221V2_7TV50

MACRO OAI222V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222V1_7TV50 0 0 ;
  SIZE 7.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.86 1.56 5.26 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.815 1.56 6.16 2 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.49 1.52 2.76 2.055 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.305 1.52 3.72 1.99 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.885 2.01 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.525 0.95 0.855 1.39 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.48 2.405 0.76 3.48 ;
        RECT 3.68 2.795 3.96 3.48 ;
        RECT 6.19 2.405 6.47 3.48 ;
        RECT 0 3.24 7.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.66 -0.12 4.94 0.565 ;
        RECT 6.46 -0.12 6.74 0.565 ;
        RECT 0 -0.12 7.2 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.17 0.71 1.36 2.525 ;
        RECT 1.12 0.71 1.41 0.9 ;
        RECT 1.17 2.335 4.87 2.525 ;
        RECT 4.4 2.335 4.72 2.76 ;
        RECT 4.4 2.335 4.87 2.53 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.625 -0.24 3.675 1.555 ;
        RECT -0.12 -0.24 7.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.625 3.94 ;
        RECT 3.675 1.46 7.78 3.94 ;
        RECT -0.58 1.555 7.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.545 0.32 4.04 0.51 ;
      RECT 0.17 0.38 0.685 0.57 ;
      RECT 2.09 0.32 2.37 0.57 ;
      RECT 3.89 0.38 4.29 0.57 ;
      RECT 3.05 0.71 3.33 0.96 ;
      RECT 5.605 0.33 5.795 0.96 ;
      RECT 3.05 0.77 5.795 0.96 ;
  END
END OAI222V1_7TV50

MACRO OAI222V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222V2_7TV50 0 0 ;
  SIZE 12.96 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.105 1.92 10.48 2.28 ;
        RECT 10.105 1.92 11.235 2.11 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.2 1.49 9.52 1.8 ;
        RECT 9.2 1.49 12.04 1.68 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8 1.96 7.12 2.28 ;
        RECT 6.395 1.96 7.585 2.15 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.59 1.56 5.78 2.2 ;
        RECT 5.59 1.56 8.56 1.75 ;
        RECT 8.235 1.56 8.56 1.8 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.99 1.56 2.32 1.8 ;
        RECT 1.99 1.61 3.13 1.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.225 1.915 1.415 2.23 ;
        RECT 2.48 2.04 2.8 2.28 ;
        RECT 3.635 1.915 3.825 2.23 ;
        RECT 1.225 2.04 3.825 2.23 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.705 2.405 0.985 3.48 ;
        RECT 4.125 2.97 4.405 3.48 ;
        RECT 8.765 2.97 9.045 3.48 ;
        RECT 12.235 2.405 12.515 3.48 ;
        RECT 0 3.24 12.96 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 9.58 -0.12 9.86 0.565 ;
        RECT 11.38 -0.12 11.66 0.565 ;
        RECT 0 -0.12 12.96 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 2.52 3.28 2.76 ;
        RECT 1.455 0.765 4.465 0.955 ;
        RECT 4.275 0.765 4.465 2.76 ;
        RECT 2.405 2.57 10.825 2.76 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.58 -0.24 7.49 1.585 ;
        RECT -0.12 -0.24 13.08 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.58 3.94 ;
        RECT 7.49 1.46 13.54 3.94 ;
        RECT -0.58 1.585 13.54 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.495 0.375 8.06 0.565 ;
      RECT 8.725 0.57 8.915 0.955 ;
      RECT 10.525 0.58 10.715 0.955 ;
      RECT 12.325 0.58 12.515 0.955 ;
      RECT 5.02 0.765 12.515 0.955 ;
  END
END OAI222V2_7TV50

MACRO OAI22BBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22BBV1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.36 1.51 1.8 1.905 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.495 1.03 1.03 1.385 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.75 1.53 4.275 1.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.67 1.56 5.2 1.875 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.305 2.37 0.585 3.48 ;
        RECT 2.535 2.79 2.815 3.48 ;
        RECT 5.045 2.4 5.325 3.48 ;
        RECT 2.535 3.235 5.325 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 -0.12 0.535 0.83 ;
        RECT 4.345 -0.12 4.625 0.58 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 0.6 2.94 0.84 ;
        RECT 2.75 0.6 2.94 2.43 ;
        RECT 2.75 2.24 3.725 2.43 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2 1.065 2.55 1.36 ;
      RECT 2 0.595 2.19 2.43 ;
      RECT 1.155 2.24 2.19 2.43 ;
      RECT 3.49 0.595 3.68 0.97 ;
      RECT 5.29 0.595 5.48 0.97 ;
      RECT 3.49 0.78 5.48 0.97 ;
  END
END OAI22BBV1_7TV50

MACRO OAI22BBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22BBV2_7TV50 0 0 ;
  SIZE 8.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.04 1.61 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.52 0.84 1.84 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8 1.08 7.12 1.32 ;
        RECT 5.825 1.125 7.12 1.32 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.875 1.55 5.2 1.8 ;
        RECT 4.875 1.6 8 1.8 ;
        RECT 7.81 1.6 8 2.04 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.2 2.405 0.48 3.48 ;
        RECT 1.9 2.405 2.18 3.48 ;
        RECT 2.49 2.405 2.77 3.48 ;
        RECT 4.41 2.795 4.69 3.48 ;
        RECT 8.14 2.4 8.42 3.48 ;
        RECT 0 3.24 8.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.66 ;
        RECT 5.31 -0.12 5.59 0.435 ;
        RECT 7.23 -0.12 7.51 0.435 ;
        RECT 0 -0.12 8.64 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.39 0.71 3.67 0.9 ;
        RECT 3.48 0.71 3.67 2.545 ;
        RECT 3.48 1.52 3.72 1.84 ;
        RECT 3.48 2.355 6.55 2.545 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.655 -0.24 4.145 1.53 ;
        RECT -0.12 -0.24 8.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.655 3.94 ;
        RECT 4.145 1.46 9.22 3.94 ;
        RECT -0.58 1.53 9.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.945 0.595 2.135 2.065 ;
      RECT 1.095 1.875 3.145 2.065 ;
      RECT 1.095 1.875 1.285 2.545 ;
      RECT 2.535 0.32 4.585 0.51 ;
      RECT 4.39 0.32 4.585 0.825 ;
      RECT 2.535 0.32 2.725 0.7 ;
      RECT 4.39 0.635 8.47 0.825 ;
  END
END OAI22BBV2_7TV50

MACRO OAI22V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.47 1.375 2.8 2.015 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.29 1.765 3.485 2.28 ;
        RECT 3.29 2.01 3.76 2.28 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.52 1.93 2.09 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.49 0.95 0.88 1.32 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.425 2.405 0.705 3.48 ;
        RECT 3.825 2.795 4.105 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.975 -0.12 3.255 0.565 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.71 1.27 2.615 ;
        RECT 1.08 2 1.32 2.615 ;
        RECT 1.08 0.71 1.395 0.9 ;
        RECT 1.08 2.425 2.305 2.615 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.58 -0.24 1.79 1.53 ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.58 3.94 ;
        RECT 1.79 1.46 4.9 3.94 ;
        RECT -0.58 1.53 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 0.32 2.31 0.51 ;
      RECT 0.2 0.32 0.39 0.61 ;
      RECT 2.12 0.32 2.31 0.955 ;
      RECT 3.92 0.58 4.11 0.955 ;
      RECT 2.12 0.765 4.11 0.955 ;
  END
END OAI22V1_7TV50

MACRO OAI22V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.865 1.04 6.12 1.425 ;
        RECT 5.28 1.225 6.12 1.425 ;
        RECT 5.28 1.235 6.62 1.425 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.65 1.76 7.24 1.95 ;
        RECT 6.84 1.76 7.24 2.32 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.545 1.995 1.825 2.32 ;
        RECT 1.545 1.995 2.785 2.185 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.515 1.52 0.955 1.84 ;
        RECT 0.515 1.52 3.535 1.71 ;
        RECT 3.345 1.52 3.535 2.16 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.365 2.405 0.645 3.48 ;
        RECT 3.785 2.775 4.065 3.48 ;
        RECT 7.375 2.625 7.655 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 4.905 -0.12 5.185 0.625 ;
        RECT 6.74 -0.12 7.02 0.645 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.125 0.72 1.405 1.055 ;
        RECT 2.04 2.385 2.3 2.8 ;
        RECT 3.045 0.72 3.325 1.055 ;
        RECT 1.125 0.855 3.925 1.055 ;
        RECT 3.735 0.855 3.925 2.575 ;
        RECT 2.04 2.385 6.055 2.575 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.58 -0.24 3.75 1.615 ;
        RECT 0.58 -0.24 7.375 1.505 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.58 3.94 ;
        RECT 3.75 1.505 8.74 3.94 ;
        RECT 7.375 1.46 8.74 3.94 ;
        RECT -0.58 1.615 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 0.32 4.53 0.51 ;
      RECT 2.085 0.32 2.365 0.605 ;
      RECT 4.005 0.32 4.53 0.605 ;
      RECT 0.2 0.32 0.39 0.61 ;
      RECT 5.475 0.59 6.53 0.78 ;
      RECT 4.34 0.32 4.53 1.015 ;
      RECT 6.34 0.59 6.53 1.035 ;
      RECT 5.475 0.59 5.665 1.015 ;
      RECT 4.34 0.825 5.665 1.015 ;
      RECT 7.68 0.56 7.875 1.035 ;
      RECT 6.34 0.845 7.875 1.035 ;
  END
END OAI22V2_7TV50

MACRO OAI22XBV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22XBV1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.93 1.52 4.2 2.11 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.835 1.52 5.16 2.045 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 1.485 3.24 2.065 ;
        RECT 3 1.875 3.315 2.065 ;
    END
  END B1
  PIN B2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.52 1.08 1.84 ;
        RECT 0.89 1.52 1.08 2.095 ;
    END
  END B2N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.41 2.32 0.69 3.48 ;
        RECT 1.91 2.405 2.19 3.48 ;
        RECT 5.165 2.405 5.445 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.465 -0.12 0.655 0.875 ;
        RECT 4.73 -0.12 5.01 0.635 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 1.52 2.76 1.84 ;
        RECT 2.57 0.71 2.76 2.5 ;
        RECT 2.57 0.71 3.09 0.9 ;
        RECT 2.57 2.31 3.79 2.5 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.575 -0.24 3.7 1.53 ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.575 3.94 ;
        RECT 3.7 1.46 6.82 3.94 ;
        RECT -0.58 1.53 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.365 1.84 2.32 2.03 ;
      RECT 2.13 1.795 2.32 2.075 ;
      RECT 1.365 0.595 1.555 2.545 ;
      RECT 1.955 0.32 4.005 0.51 ;
      RECT 3.815 0.32 4.005 1.025 ;
      RECT 1.955 0.32 2.145 0.945 ;
      RECT 5.735 0.59 5.925 1.025 ;
      RECT 3.815 0.835 5.925 1.025 ;
  END
END OAI22XBV1_7TV50

MACRO OAI22XBV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22XBV2_7TV50 0 0 ;
  SIZE 10.08 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.16 1.59 8.56 1.78 ;
        RECT 8.24 1.56 8.56 1.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8 1.07 7.12 1.32 ;
        RECT 6.165 1.07 9.375 1.26 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.56 3.76 1.8 ;
        RECT 3.355 1.58 4.595 1.77 ;
    END
  END B1
  PIN B2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.02 1.04 1.32 ;
    END
  END B2N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.465 2.61 0.745 3.48 ;
        RECT 1.97 2.795 2.25 3.48 ;
        RECT 5.69 2.795 5.97 3.48 ;
        RECT 9.315 2.405 9.595 3.48 ;
        RECT 0 3.24 10.08 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.415 -0.12 0.695 0.73 ;
        RECT 6.65 -0.12 6.93 0.435 ;
        RECT 8.57 -0.12 8.85 0.435 ;
        RECT 0 -0.12 10.08 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.93 0.74 3.21 1.125 ;
        RECT 4.73 0.74 5.01 1.125 ;
        RECT 2.93 0.935 5.01 1.125 ;
        RECT 4.76 1.08 5.79 1.27 ;
        RECT 5.36 1.08 5.79 1.32 ;
        RECT 5.6 1.08 5.79 2.595 ;
        RECT 3.875 2.405 7.84 2.595 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.39 -0.24 5.55 1.56 ;
        RECT -0.12 -0.24 10.2 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.39 3.94 ;
        RECT 5.55 1.46 10.66 3.94 ;
        RECT -0.58 1.56 10.66 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.36 1.905 3 2.095 ;
      RECT 5.21 1.86 5.4 2.19 ;
      RECT 2.81 2 5.4 2.19 ;
      RECT 1.36 0.585 1.55 2.475 ;
      RECT 1.97 0.35 5.925 0.54 ;
      RECT 5.735 0.35 5.925 0.825 ;
      RECT 1.97 0.35 2.25 0.715 ;
      RECT 3.83 0.35 4.11 0.735 ;
      RECT 5.735 0.635 9.81 0.825 ;
  END
END OAI22XBV2_7TV50

MACRO OAI2XB11V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB11V1_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.39 1.56 3.81 1.905 ;
    END
  END A1
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 1.08 1.36 ;
    END
  END A2N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.25 1.52 4.73 1.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.15 1.04 5.64 1.36 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.41 2.25 0.69 3.48 ;
        RECT 1.91 2.4 2.19 3.48 ;
        RECT 4.63 2.79 4.91 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.35 -0.12 0.63 0.83 ;
        RECT 2.87 -0.12 3.15 0.64 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.53 0.5 6.07 0.69 ;
        RECT 5.88 0.5 6.07 2.43 ;
        RECT 3.78 2.24 6.07 2.43 ;
        RECT 5.88 1.52 6.12 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.365 1.805 2.64 1.995 ;
      RECT 1.365 0.595 1.555 2.475 ;
      RECT 1.955 0.59 2.145 1.03 ;
      RECT 3.875 0.59 4.065 1.03 ;
      RECT 1.955 0.84 4.065 1.03 ;
  END
END OAI2XB11V1_7TV50

MACRO OAI2XB11V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB11V2_7TV50 0 0 ;
  SIZE 9.6 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.56 3.76 1.8 ;
        RECT 3.11 1.56 4.24 1.75 ;
    END
  END A1
  PIN A2N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.395 1.02 0.88 1.32 ;
    END
  END A2N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.73 1.56 6.16 1.8 ;
        RECT 5.73 1.61 8.635 1.8 ;
        RECT 8.445 1.565 8.635 1.845 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.36 1.04 6.605 1.395 ;
        RECT 6.36 1.15 6.81 1.395 ;
        RECT 6.36 1.205 7.855 1.395 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.215 2.615 0.495 3.48 ;
        RECT 1.735 2.405 2.015 3.48 ;
        RECT 5.245 2.83 5.525 3.48 ;
        RECT 7.115 2.83 7.395 3.48 ;
        RECT 8.935 2.83 9.215 3.48 ;
        RECT 0 3.24 9.6 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.12 0.445 0.705 ;
        RECT 2.635 -0.12 2.915 0.635 ;
        RECT 4.455 -0.12 4.735 0.635 ;
        RECT 0 -0.12 9.6 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.115 0.72 7.395 0.955 ;
        RECT 7.115 0.765 8.43 0.955 ;
        RECT 8.24 0.765 8.43 1.33 ;
        RECT 8.24 1.08 8.56 1.33 ;
        RECT 8.24 1.14 9.025 1.33 ;
        RECT 8.835 1.14 9.025 2.63 ;
        RECT 3.585 2.44 9.025 2.63 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 6.41 -0.24 7.88 1.54 ;
        RECT -0.12 -0.24 9.72 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.41 3.94 ;
        RECT 7.88 1.46 10.18 3.94 ;
        RECT -0.58 1.54 10.18 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.11 1.765 2.345 1.955 ;
      RECT 2.155 1.765 2.345 2.19 ;
      RECT 4.855 1.765 5.045 2.19 ;
      RECT 2.155 2 5.045 2.19 ;
      RECT 1.11 0.54 1.3 2.48 ;
      RECT 5.4 0.325 9.155 0.515 ;
      RECT 8.875 0.325 9.155 0.635 ;
      RECT 1.78 0.595 1.97 1.025 ;
      RECT 3.58 0.595 3.77 1.025 ;
      RECT 5.4 0.325 5.59 1.025 ;
      RECT 1.78 0.835 5.59 1.025 ;
  END
END OAI2XB11V2_7TV50

MACRO OAI2XB1V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.91 1.56 4.52 1.8 ;
        RECT 4.24 1.56 4.52 1.935 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.95 1.56 3.285 1.935 ;
        RECT 2.95 1.745 3.605 1.935 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.435 1.515 0.905 1.86 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.235 2.25 0.515 3.48 ;
        RECT 1.98 2.4 2.26 3.48 ;
        RECT 4.7 2.79 4.98 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.185 -0.12 0.465 0.83 ;
        RECT 2.89 -0.12 3.17 0.64 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.75 0.64 5.11 0.83 ;
        RECT 4.92 0.64 5.11 2.43 ;
        RECT 3.85 2.24 5.11 2.43 ;
        RECT 4.92 1.52 5.16 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.385 1.805 2.665 1.995 ;
      RECT 1.385 0.595 1.575 2.475 ;
      RECT 1.975 0.59 2.165 1.03 ;
      RECT 3.895 0.59 4.085 1.03 ;
      RECT 1.975 0.84 4.085 1.03 ;
  END
END OAI2XB1V1_7TV50

MACRO OAI2XB1V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2XB1V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.8 1.83 7.345 2.285 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.25 1.48 3.44 1.8 ;
        RECT 3.25 1.56 3.76 1.8 ;
        RECT 3.25 1.61 4.285 1.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.42 1 0.88 1.32 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.305 2.61 0.585 3.48 ;
        RECT 1.88 2.405 2.16 3.48 ;
        RECT 5.43 2.795 5.71 3.48 ;
        RECT 7.165 2.795 7.445 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 -0.12 0.535 0.765 ;
        RECT 2.73 -0.12 3.01 0.635 ;
        RECT 4.53 -0.12 4.81 0.635 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.36 0.71 6.55 2.595 ;
        RECT 6.36 1.52 6.6 1.84 ;
        RECT 3.58 2.405 6.6 2.595 ;
        RECT 6.36 0.71 6.67 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 5.96 -0.24 7.545 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.96 3.94 ;
        RECT 7.545 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.2 1.81 2.57 2 ;
      RECT 4.95 1.765 5.14 2.19 ;
      RECT 2.38 2 5.14 2.19 ;
      RECT 1.2 0.565 1.39 2.475 ;
      RECT 5.475 0.32 7.585 0.51 ;
      RECT 7.395 0.32 7.585 0.685 ;
      RECT 1.875 0.595 2.065 1.025 ;
      RECT 3.675 0.595 3.865 1.025 ;
      RECT 5.475 0.32 5.665 1.025 ;
      RECT 1.875 0.835 5.665 1.025 ;
  END
END OAI2XB1V2_7TV50

MACRO OAI31V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 1.56 2.81 2.055 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4 1.805 1.87 2.32 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.485 1.475 0.955 1.99 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.34 1.01 3.72 1.495 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 2.4 0.445 3.48 ;
        RECT 3.565 2.79 3.845 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.165 -0.12 0.445 0.58 ;
        RECT 1.965 -0.12 2.245 0.58 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.765 0.605 4.11 0.795 ;
        RECT 3.92 0.605 4.11 2.445 ;
        RECT 2.715 2.255 4.11 2.445 ;
        RECT 3.92 1.52 4.2 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.11 0.595 1.3 0.97 ;
      RECT 2.91 0.595 3.1 0.97 ;
      RECT 1.11 0.78 3.1 0.97 ;
  END
END OAI31V1_7TV50

MACRO OAI31V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31V2_7TV50 0 0 ;
  SIZE 8.64 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.48 2.035 2.83 2.28 ;
        RECT 2.48 2.035 3.8 2.225 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2 1.56 2.32 1.8 ;
        RECT 1.55 1.61 4.7 1.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.08 1.84 1.32 ;
        RECT 0.765 1.125 5.45 1.315 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.295 1.505 7.745 1.84 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.405 0.435 3.48 ;
        RECT 5.7 2.795 5.98 3.48 ;
        RECT 7.625 2.405 7.905 3.48 ;
        RECT 0 3.24 8.64 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.115 -0.12 1.395 0.435 ;
        RECT 3.035 -0.12 3.315 0.435 ;
        RECT 4.955 -0.12 5.235 0.435 ;
        RECT 0 -0.12 8.64 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.085 2.57 4.405 2.76 ;
        RECT 6.36 1.52 6.6 1.84 ;
        RECT 6.41 0.71 6.6 2.595 ;
        RECT 4.215 2.405 7.055 2.595 ;
        RECT 6.41 0.71 7.145 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.07 -0.24 8.06 1.53 ;
        RECT -0.12 -0.24 8.76 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.07 3.94 ;
        RECT 8.06 1.46 9.22 3.94 ;
        RECT -0.58 1.53 9.22 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 5.96 0.32 8.06 0.51 ;
      RECT 7.87 0.32 8.06 0.615 ;
      RECT 5.96 0.32 6.15 0.825 ;
      RECT 0.155 0.635 6.15 0.825 ;
  END
END OAI31V2_7TV50

MACRO OAI32V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32V1_7TV50 0 0 ;
  SIZE 5.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.495 1.52 2.86 1.99 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.55 1.44 1.91 1.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.97 1.62 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.38 1.52 3.76 1.99 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.405 1.52 4.805 1.99 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.265 2.405 0.545 3.48 ;
        RECT 4.72 2.405 5 3.48 ;
        RECT 0 3.24 5.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.265 -0.12 0.545 0.565 ;
        RECT 2.065 -0.12 2.345 0.565 ;
        RECT 0 -0.12 5.76 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 0.71 4.2 1.36 ;
        RECT 4.01 0.71 4.2 2.595 ;
        RECT 3 2.405 4.2 2.595 ;
        RECT 3.91 0.71 4.205 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 3.495 -0.24 5.18 1.53 ;
        RECT -0.12 -0.24 5.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.495 3.94 ;
        RECT 5.18 1.46 6.34 3.94 ;
        RECT -0.58 1.53 6.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 3.01 0.32 5.12 0.51 ;
      RECT 4.93 0.32 5.12 0.63 ;
      RECT 1.21 0.58 1.4 0.955 ;
      RECT 3.01 0.32 3.2 0.955 ;
      RECT 1.21 0.765 3.2 0.955 ;
  END
END OAI32V1_7TV50

MACRO OAI32V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32V2_7TV50 0 0 ;
  SIZE 10.56 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.81 1.875 3.28 2.28 ;
        RECT 2.81 1.875 4.16 2.065 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.045 1.39 5.16 1.58 ;
        RECT 4.8 1.39 5.16 1.84 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.035 0.98 1.36 1.32 ;
        RECT 1.035 0.98 6.015 1.18 ;
        RECT 5.825 0.98 6.015 1.37 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.67 1.875 8.08 2.28 ;
        RECT 7.67 1.875 8.945 2.065 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.84 1.04 7.035 1.84 ;
        RECT 6.84 1.21 7.08 1.84 ;
        RECT 6.84 1.21 9.88 1.4 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.515 2.395 0.795 3.48 ;
        RECT 6.095 2.97 6.375 3.48 ;
        RECT 10.06 2.795 10.34 3.48 ;
        RECT 0 3.24 10.56 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.475 -0.12 1.755 0.39 ;
        RECT 3.395 -0.12 3.675 0.39 ;
        RECT 5.315 -0.12 5.595 0.39 ;
        RECT 0 -0.12 10.56 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.235 0.71 7.515 1.01 ;
        RECT 9.115 2.36 9.305 2.77 ;
        RECT 3.505 2.58 9.305 2.77 ;
        RECT 9.155 0.71 9.435 1.01 ;
        RECT 7.235 0.82 10.27 1.01 ;
        RECT 10.08 0.82 10.27 2.55 ;
        RECT 9.115 2.36 10.27 2.55 ;
        RECT 10.08 1.52 10.44 1.84 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 5.91 -0.24 9.98 1.53 ;
        RECT -0.12 -0.24 10.68 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.91 3.94 ;
        RECT 9.98 1.46 11.14 3.94 ;
        RECT -0.58 1.53 11.14 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 6.345 0.32 10.35 0.51 ;
      RECT 8.24 0.32 8.43 0.62 ;
      RECT 10.16 0.32 10.35 0.62 ;
      RECT 6.345 0.32 6.555 0.78 ;
      RECT 0.515 0.59 6.555 0.78 ;
  END
END OAI32V2_7TV50

MACRO OR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2V1_7TV50 0 0 ;
  SIZE 3.36 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.41 1.04 0.87 1.36 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.52 1.56 1.93 1.915 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.065 2.79 2.345 3.48 ;
        RECT 0 3.24 3.36 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.2 -0.12 0.48 0.83 ;
        RECT 2.015 -0.12 2.295 0.83 ;
        RECT 0 -0.12 3.36 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.96 0.595 3.15 2.475 ;
        RECT 2.96 1.04 3.24 1.36 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 3.48 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.94 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.115 0.64 1.395 0.83 ;
      RECT 1.115 0.64 1.315 2.43 ;
      RECT 1.115 2.23 2.675 2.43 ;
      RECT 2.485 1.76 2.675 2.43 ;
      RECT 0.365 2.24 2.675 2.43 ;
  END
END OR2V1_7TV50

MACRO OR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2V2_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.47 1.56 0.95 1.86 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.55 1.04 1.97 1.385 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.05 2.66 2.33 3.48 ;
        RECT 3.85 2.4 4.13 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.25 -0.12 0.53 0.66 ;
        RECT 2.05 -0.12 2.33 0.66 ;
        RECT 3.85 -0.12 4.13 0.58 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3 0.555 3.19 2.475 ;
        RECT 2.95 0.555 3.24 0.745 ;
        RECT 3 1.52 3.24 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.15 0.555 1.43 0.745 ;
      RECT 1.15 0.555 1.35 2.43 ;
      RECT 1.15 2.23 2.66 2.43 ;
      RECT 2.47 1.76 2.66 2.43 ;
      RECT 0.28 2.24 2.66 2.43 ;
  END
END OR2V2_7TV50

MACRO OR2V4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2V4_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.81 1.8 2.32 ;
        RECT 1.56 1.81 2.945 2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.065 1.42 3.76 1.61 ;
        RECT 3.43 1.42 3.76 1.8 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.49 2.555 0.77 3.48 ;
        RECT 3.965 2.81 4.245 3.48 ;
        RECT 5.79 2.405 6.07 3.48 ;
        RECT 7.64 2.405 7.92 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.44 -0.12 0.72 0.73 ;
        RECT 2.24 -0.12 2.52 0.73 ;
        RECT 4.04 -0.12 4.32 0.73 ;
        RECT 5.84 -0.12 6.12 0.565 ;
        RECT 7.64 -0.12 7.92 0.565 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.92 1.04 5.175 1.36 ;
        RECT 4.985 0.595 5.175 2.48 ;
        RECT 4.985 1.21 6.975 1.4 ;
        RECT 6.785 0.595 6.975 2.48 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.385 0.595 1.575 1.12 ;
      RECT 3.185 0.595 3.375 1.12 ;
      RECT 1.385 0.93 4.695 1.12 ;
      RECT 4.505 0.93 4.695 2.435 ;
      RECT 2.29 2.245 4.695 2.435 ;
  END
END OR2V4_7TV50

MACRO OR3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3V1_7TV50 0 0 ;
  SIZE 4.32 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.945 1.575 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.515 1.56 1.84 2.005 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.445 1.42 2.805 1.835 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.035 2.4 3.315 3.48 ;
        RECT 0 3.24 4.32 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 -0.12 1.405 0.44 ;
        RECT 2.985 -0.12 3.265 0.83 ;
        RECT 0 -0.12 4.32 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.93 0.595 4.2 0.875 ;
        RECT 3.96 1.52 4.2 1.84 ;
        RECT 4.01 0.595 4.2 2.475 ;
        RECT 3.93 2.195 4.2 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 4.44 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.9 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.165 0.64 2.505 0.83 ;
      RECT 2.315 0.64 2.505 1.22 ;
      RECT 2.315 1.03 3.595 1.22 ;
      RECT 3.405 1.03 3.595 1.31 ;
      RECT 0.165 0.64 0.355 2.43 ;
      RECT 0.165 2.24 0.615 2.43 ;
  END
END OR3V1_7TV50

MACRO OR3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3V2_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.76 0.845 2.32 ;
        RECT 0.6 1.76 0.875 2.04 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.555 1.76 1.8 2.32 ;
        RECT 1.555 1.76 1.83 2.04 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.4 1.435 2.8 1.8 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 2.815 2.27 3.095 3.48 ;
        RECT 4.665 2.4 4.945 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 -0.12 1.345 0.66 ;
        RECT 2.865 -0.12 3.145 0.66 ;
        RECT 4.665 -0.12 4.945 0.58 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.765 0.64 4.15 0.83 ;
        RECT 3.96 0.64 4.15 2.475 ;
        RECT 3.805 2.285 4.15 2.475 ;
        RECT 3.96 1.52 4.2 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.01 0.595 2.2 1.22 ;
      RECT 0.21 1.02 2.2 1.22 ;
      RECT 0.21 1.03 3.49 1.22 ;
      RECT 3.3 1.03 3.49 1.31 ;
      RECT 0.21 0.595 0.4 2.475 ;
  END
END OR3V2_7TV50

MACRO OR4V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.56 1.56 1.07 1.845 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.46 1.465 1.84 1.895 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.65 1.52 3.24 1.895 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.465 3.72 1.98 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.98 2.4 4.26 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.33 -0.12 0.61 0.83 ;
        RECT 2.13 -0.12 2.41 0.83 ;
        RECT 3.93 -0.12 4.21 0.83 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.875 0.595 5.065 2.475 ;
        RECT 4.875 1.52 5.16 1.84 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.275 0.595 1.465 1.265 ;
      RECT 3.075 0.595 3.265 1.265 ;
      RECT 1.275 1.075 4.635 1.265 ;
      RECT 2.04 1.075 2.23 2.43 ;
      RECT 0.38 2.24 2.23 2.43 ;
  END
END OR4V1_7TV50

MACRO OR4V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4V2_7TV50 0 0 ;
  SIZE 6.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.76 1.34 2.33 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 1.415 1.9 1.84 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.5 1.805 2.83 2.33 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.445 1.47 3.855 1.95 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 3.84 2.27 4.12 3.48 ;
        RECT 5.775 2.4 6.055 3.48 ;
        RECT 0 3.24 6.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.375 -0.12 0.655 0.58 ;
        RECT 2.175 -0.12 2.455 0.58 ;
        RECT 3.975 -0.12 4.255 0.58 ;
        RECT 5.775 -0.12 6.055 0.58 ;
        RECT 0 -0.12 6.24 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.92 0.46 5.11 2.475 ;
        RECT 4.92 0.56 5.16 0.88 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 6.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 6.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.32 0.595 1.51 1 ;
      RECT 3.12 0.595 3.31 1 ;
      RECT 0.65 0.81 4.585 1 ;
      RECT 4.395 0.81 4.585 1.31 ;
      RECT 0.65 0.81 0.84 2.475 ;
  END
END OR4V2_7TV50

MACRO PULL0_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN PULL0_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.08 2.38 1.36 3.48 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.18 -0.12 0.46 0.79 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.505 1.44 0.905 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.265 1.945 0.475 2.66 ;
  END
END PULL0_7TV50

MACRO PULL1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN PULL1_7TV50 0 0 ;
  SIZE 1.92 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.4 2.275 0.68 3.48 ;
        RECT 0 3.24 1.92 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.3 -0.12 1.58 0.86 ;
        RECT 0 -0.12 1.92 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 2.04 1.53 2.28 ;
        RECT 1.25 2.04 1.53 2.43 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.04 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.5 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.435 0.595 0.645 1.31 ;
  END
END PULL1_7TV50

MACRO SDQNV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDQNV1_7TV50 0 0 ;
  SIZE 16.8 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.76 1.56 6.36 1.8 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.945 2.41 2.335 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.11 0.56 16.3 2.48 ;
        RECT 16.11 0.56 16.68 0.88 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.265 ;
        RECT 0.6 1.075 3.41 1.265 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.08 1.605 4.68 1.84 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.605 1.285 3.48 ;
        RECT 4.265 2.97 4.545 3.48 ;
        RECT 9.965 2.44 10.245 3.48 ;
        RECT 13.39 2.44 13.67 3.48 ;
        RECT 15.215 2.28 15.495 3.48 ;
        RECT 0 3.24 16.8 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.875 ;
        RECT 4.455 -0.12 4.69 0.875 ;
        RECT 6.135 -0.12 6.415 0.97 ;
        RECT 10.285 -0.12 10.565 0.555 ;
        RECT 13.905 -0.12 14.185 0.82 ;
        RECT 15.395 -0.12 15.675 0.625 ;
        RECT 0 -0.12 16.8 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.83 -0.24 7.72 1.6 ;
        RECT 4.83 -0.24 11.83 1.53 ;
        RECT -0.12 -0.24 16.92 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.83 3.94 ;
        RECT 7.72 1.53 17.38 3.94 ;
        RECT 11.83 1.46 17.38 3.94 ;
        RECT -0.58 1.6 17.38 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.485 3.215 1.675 ;
      RECT 3.025 1.485 3.215 2.37 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.28 2.025 6.65 2.215 ;
      RECT 5.28 0.735 5.47 2.65 ;
      RECT 5.19 2.46 5.47 2.65 ;
      RECT 2.605 2.575 4.935 2.765 ;
      RECT 4.745 2.575 4.935 3.04 ;
      RECT 7.56 2.52 7.75 3.04 ;
      RECT 4.745 2.85 7.75 3.04 ;
      RECT 4.89 0.345 5.935 0.535 ;
      RECT 2.755 0.64 3.875 0.83 ;
      RECT 7.625 0.71 7.905 0.9 ;
      RECT 3.685 0.64 3.875 1.265 ;
      RECT 5.745 0.345 5.935 1.36 ;
      RECT 4.89 0.345 5.08 1.265 ;
      RECT 3.685 1.075 5.08 1.265 ;
      RECT 7.625 0.71 7.815 1.36 ;
      RECT 5.745 1.17 7.815 1.36 ;
      RECT 8.495 0.71 8.805 0.9 ;
      RECT 8.495 1.535 10.62 1.725 ;
      RECT 8.495 0.71 8.685 2.595 ;
      RECT 8.365 2.405 8.685 2.595 ;
      RECT 8.885 1.925 11.245 2.115 ;
      RECT 8.885 1.925 9.075 2.205 ;
      RECT 11.055 1.925 11.245 2.205 ;
      RECT 11.245 0.71 11.635 0.9 ;
      RECT 9.7 1.145 11.635 1.335 ;
      RECT 11.445 0.71 11.635 2.595 ;
      RECT 10.815 2.405 11.635 2.595 ;
      RECT 7.125 0.32 9.33 0.51 ;
      RECT 10.83 0.32 12.05 0.51 ;
      RECT 10.83 0.32 11.02 0.945 ;
      RECT 9.14 0.755 11.02 0.945 ;
      RECT 7.125 0.32 7.315 0.97 ;
      RECT 7.035 0.78 7.315 0.97 ;
      RECT 9.14 0.32 9.33 1.335 ;
      RECT 9.05 1.145 9.33 1.335 ;
      RECT 11.86 0.32 12.05 2.16 ;
      RECT 8.105 0.32 8.295 2.16 ;
      RECT 6.935 1.97 8.295 2.16 ;
      RECT 11.86 1.97 12.445 2.16 ;
      RECT 6.935 1.97 7.125 2.65 ;
      RECT 6.845 2.46 7.125 2.65 ;
      RECT 12.25 0.54 12.44 0.82 ;
      RECT 12.25 0.63 12.835 0.82 ;
      RECT 12.645 1.81 14.21 2 ;
      RECT 12.645 0.63 12.835 2.59 ;
      RECT 11.835 2.4 12.835 2.59 ;
      RECT 11.835 2.4 12.025 2.68 ;
      RECT 14.54 0.345 14.73 1.21 ;
      RECT 13.53 1.02 14.73 1.21 ;
      RECT 14.41 1.02 14.6 2.48 ;
  END
END SDQNV1_7TV50

MACRO SDQNV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDQNV2_7TV50 0 0 ;
  SIZE 17.76 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.76 1.56 6.36 1.8 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.945 2.41 2.335 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.11 0.56 16.3 2.48 ;
        RECT 16.11 0.56 16.68 0.88 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.265 ;
        RECT 0.6 1.075 3.41 1.265 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.08 1.605 4.68 1.84 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.51 1.285 3.48 ;
        RECT 4.265 2.97 4.545 3.48 ;
        RECT 9.965 2.44 10.245 3.48 ;
        RECT 13.39 2.62 13.67 3.48 ;
        RECT 15.215 2.28 15.495 3.48 ;
        RECT 16.92 2.28 17.2 3.48 ;
        RECT 0 3.24 17.76 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.84 ;
        RECT 4.455 -0.12 4.69 0.805 ;
        RECT 6.135 -0.12 6.415 0.97 ;
        RECT 10.285 -0.12 10.565 0.555 ;
        RECT 13.905 -0.12 14.185 0.82 ;
        RECT 15.395 -0.12 15.675 0.625 ;
        RECT 17.195 -0.12 17.475 0.725 ;
        RECT 0 -0.12 17.76 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.83 -0.24 7.72 1.6 ;
        RECT 4.83 -0.24 11.83 1.53 ;
        RECT -0.12 -0.24 17.88 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.83 3.94 ;
        RECT 7.72 1.53 18.34 3.94 ;
        RECT 11.83 1.46 18.34 3.94 ;
        RECT -0.58 1.6 18.34 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.485 3.215 1.675 ;
      RECT 3.025 1.485 3.215 2.18 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.28 2.025 6.65 2.215 ;
      RECT 5.28 0.735 5.47 2.65 ;
      RECT 5.19 2.46 5.47 2.65 ;
      RECT 2.605 2.575 4.935 2.765 ;
      RECT 4.745 2.575 4.935 3.04 ;
      RECT 7.56 2.64 7.75 3.04 ;
      RECT 4.745 2.85 7.75 3.04 ;
      RECT 4.89 0.345 5.935 0.535 ;
      RECT 2.755 0.57 3.875 0.76 ;
      RECT 7.625 0.71 7.905 0.9 ;
      RECT 3.685 0.57 3.875 1.195 ;
      RECT 5.745 0.345 5.935 1.36 ;
      RECT 4.89 0.345 5.08 1.195 ;
      RECT 3.685 1.005 5.08 1.195 ;
      RECT 7.625 0.71 7.815 1.36 ;
      RECT 5.745 1.17 7.815 1.36 ;
      RECT 8.495 0.71 8.805 0.9 ;
      RECT 8.495 1.535 10.62 1.725 ;
      RECT 8.495 0.71 8.685 2.595 ;
      RECT 8.365 2.405 8.685 2.595 ;
      RECT 11.055 1.875 11.245 2.155 ;
      RECT 8.885 1.925 11.245 2.155 ;
      RECT 8.885 1.925 9.075 2.205 ;
      RECT 11.245 0.71 11.635 0.9 ;
      RECT 9.7 1.145 11.635 1.335 ;
      RECT 11.445 0.71 11.635 2.595 ;
      RECT 10.815 2.405 11.635 2.595 ;
      RECT 7.125 0.32 9.33 0.51 ;
      RECT 10.83 0.32 12.05 0.51 ;
      RECT 10.83 0.32 11.02 0.945 ;
      RECT 9.14 0.755 11.02 0.945 ;
      RECT 7.125 0.32 7.315 0.97 ;
      RECT 7.035 0.78 7.315 0.97 ;
      RECT 9.14 0.32 9.33 1.335 ;
      RECT 9.05 1.145 9.33 1.335 ;
      RECT 11.86 0.32 12.05 2.34 ;
      RECT 8.105 0.32 8.295 2.16 ;
      RECT 6.935 1.97 8.295 2.16 ;
      RECT 11.86 2.15 12.445 2.34 ;
      RECT 6.935 1.97 7.125 2.65 ;
      RECT 6.845 2.46 7.125 2.65 ;
      RECT 12.25 0.54 12.44 0.82 ;
      RECT 12.25 0.63 12.835 0.82 ;
      RECT 12.645 1.81 14.21 2 ;
      RECT 12.645 0.63 12.835 2.73 ;
      RECT 11.835 2.54 12.835 2.73 ;
      RECT 11.835 2.54 12.025 2.82 ;
      RECT 14.54 0.345 14.73 1.21 ;
      RECT 13.53 1.02 14.73 1.21 ;
      RECT 14.41 1.02 14.6 2.48 ;
  END
END SDQNV2_7TV50

MACRO SDQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDQV1_7TV50 0 0 ;
  SIZE 18.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.76 1.56 6.36 1.8 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.945 2.41 2.335 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 17.675 0.56 17.865 2.48 ;
        RECT 17.675 0.56 18.12 0.88 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.265 ;
        RECT 0.6 1.075 3.41 1.265 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.08 1.605 4.68 1.84 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.51 1.285 3.48 ;
        RECT 4.265 2.97 4.545 3.48 ;
        RECT 10.035 2.44 10.27 3.48 ;
        RECT 12.14 2.265 12.42 3.48 ;
        RECT 15.34 2.61 15.62 3.48 ;
        RECT 16.78 2.295 17.06 3.48 ;
        RECT 0 3.24 18.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.815 ;
        RECT 4.455 -0.12 4.69 0.755 ;
        RECT 6.135 -0.12 6.415 0.97 ;
        RECT 10.285 -0.12 10.565 0.555 ;
        RECT 12.115 -0.12 12.35 0.735 ;
        RECT 15.47 -0.12 15.75 0.82 ;
        RECT 16.96 -0.12 17.24 0.625 ;
        RECT 0 -0.12 18.72 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.83 -0.24 7.72 1.6 ;
        RECT 4.83 -0.24 11.83 1.53 ;
        RECT -0.12 -0.24 18.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.83 3.94 ;
        RECT 7.72 1.53 19.3 3.94 ;
        RECT 11.83 1.46 19.3 3.94 ;
        RECT -0.58 1.6 19.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.485 3.215 1.675 ;
      RECT 3.025 1.485 3.215 2.18 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.28 2.025 6.65 2.215 ;
      RECT 5.28 0.735 5.47 2.65 ;
      RECT 5.19 2.46 5.47 2.65 ;
      RECT 2.605 2.575 4.935 2.765 ;
      RECT 4.745 2.575 4.935 3.04 ;
      RECT 7.63 2.64 7.82 3.04 ;
      RECT 4.745 2.85 7.82 3.04 ;
      RECT 4.89 0.345 5.935 0.535 ;
      RECT 2.755 0.56 3.875 0.75 ;
      RECT 7.625 0.71 7.905 0.9 ;
      RECT 3.685 0.56 3.875 1.145 ;
      RECT 4.89 0.345 5.08 1.145 ;
      RECT 3.685 0.955 5.08 1.145 ;
      RECT 5.745 0.345 5.935 1.36 ;
      RECT 7.625 0.71 7.815 1.36 ;
      RECT 5.745 1.17 7.815 1.36 ;
      RECT 8.525 0.71 8.805 0.9 ;
      RECT 8.525 1.535 11 1.725 ;
      RECT 8.525 0.71 8.715 2.595 ;
      RECT 8.435 2.405 8.715 2.595 ;
      RECT 11.245 0.71 11.525 0.9 ;
      RECT 9.85 1.145 11.435 1.335 ;
      RECT 11.245 1.43 12.795 1.62 ;
      RECT 11.245 0.71 11.435 2.595 ;
      RECT 10.885 2.405 11.435 2.595 ;
      RECT 11.635 1.82 13.545 2.01 ;
      RECT 8.955 1.925 9.145 2.205 ;
      RECT 8.955 2.015 10.685 2.205 ;
      RECT 10.495 2.015 10.685 2.985 ;
      RECT 11.635 1.82 11.825 2.985 ;
      RECT 10.495 2.795 11.825 2.985 ;
      RECT 7.125 0.32 9.33 0.51 ;
      RECT 10.83 0.32 11.915 0.51 ;
      RECT 10.83 0.32 11.02 0.945 ;
      RECT 9.14 0.755 11.02 0.945 ;
      RECT 7.125 0.32 7.315 0.97 ;
      RECT 7.035 0.78 7.315 0.97 ;
      RECT 11.725 0.32 11.915 1.21 ;
      RECT 11.725 1.02 14.35 1.21 ;
      RECT 9.14 0.32 9.33 1.335 ;
      RECT 9.05 1.145 9.33 1.335 ;
      RECT 8.105 0.32 8.295 2.16 ;
      RECT 6.935 1.97 8.295 2.16 ;
      RECT 14.16 1.02 14.35 2.375 ;
      RECT 6.935 1.97 7.125 2.65 ;
      RECT 6.845 2.46 7.125 2.65 ;
      RECT 13.77 0.585 14.765 0.775 ;
      RECT 14.575 1.81 15.775 2 ;
      RECT 14.575 0.585 14.765 2.765 ;
      RECT 13.74 2.575 14.765 2.765 ;
      RECT 16.105 0.345 16.295 1.21 ;
      RECT 15.095 1.02 16.295 1.21 ;
      RECT 15.975 1.02 16.165 2.48 ;
  END
END SDQV1_7TV50

MACRO SDQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDQV2_7TV50 0 0 ;
  SIZE 19.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.76 1.56 6.36 1.8 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.945 2.41 2.335 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 17.675 0.56 17.865 2.48 ;
        RECT 17.675 0.56 18.12 0.88 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.265 ;
        RECT 0.6 1.075 3.41 1.265 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.08 1.605 4.68 1.84 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.515 1.285 3.48 ;
        RECT 4.265 2.97 4.545 3.48 ;
        RECT 10.035 2.44 10.27 3.48 ;
        RECT 12.14 2.265 12.42 3.48 ;
        RECT 15.34 2.61 15.62 3.48 ;
        RECT 16.78 2.295 17.06 3.48 ;
        RECT 18.48 2.28 18.76 3.48 ;
        RECT 0 3.24 19.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.815 ;
        RECT 4.455 -0.12 4.69 0.755 ;
        RECT 6.135 -0.12 6.415 0.97 ;
        RECT 10.285 -0.12 10.565 0.555 ;
        RECT 12.115 -0.12 12.35 0.735 ;
        RECT 15.47 -0.12 15.75 0.82 ;
        RECT 16.96 -0.12 17.24 0.625 ;
        RECT 18.76 -0.12 19.04 0.75 ;
        RECT 0 -0.12 19.2 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.83 -0.24 7.72 1.6 ;
        RECT 4.83 -0.24 11.83 1.53 ;
        RECT -0.12 -0.24 19.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.83 3.94 ;
        RECT 7.72 1.53 19.78 3.94 ;
        RECT 11.83 1.46 19.78 3.94 ;
        RECT -0.58 1.6 19.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.485 3.215 1.675 ;
      RECT 3.025 1.485 3.215 2.18 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.28 2.025 6.65 2.215 ;
      RECT 5.28 0.735 5.47 2.65 ;
      RECT 5.19 2.46 5.47 2.65 ;
      RECT 2.605 2.575 4.935 2.765 ;
      RECT 4.745 2.575 4.935 3.04 ;
      RECT 7.63 2.64 7.82 3.04 ;
      RECT 4.745 2.85 7.82 3.04 ;
      RECT 4.89 0.345 5.935 0.535 ;
      RECT 2.755 0.56 3.875 0.75 ;
      RECT 7.625 0.71 7.905 0.9 ;
      RECT 3.685 0.56 3.875 1.145 ;
      RECT 4.89 0.345 5.08 1.145 ;
      RECT 3.685 0.955 5.08 1.145 ;
      RECT 5.745 0.345 5.935 1.36 ;
      RECT 7.625 0.71 7.815 1.36 ;
      RECT 5.745 1.17 7.815 1.36 ;
      RECT 8.525 0.71 8.805 0.9 ;
      RECT 8.525 1.535 11 1.725 ;
      RECT 8.525 0.71 8.715 2.595 ;
      RECT 8.435 2.405 8.715 2.595 ;
      RECT 11.245 0.71 11.525 0.9 ;
      RECT 9.85 1.145 11.435 1.335 ;
      RECT 11.245 1.43 12.795 1.62 ;
      RECT 11.245 0.71 11.435 2.595 ;
      RECT 10.885 2.405 11.435 2.595 ;
      RECT 11.635 1.82 13.545 2.01 ;
      RECT 8.955 1.925 9.145 2.205 ;
      RECT 8.955 2.015 10.685 2.205 ;
      RECT 10.495 2.015 10.685 2.985 ;
      RECT 11.635 1.82 11.825 2.985 ;
      RECT 10.495 2.795 11.825 2.985 ;
      RECT 7.125 0.32 9.33 0.51 ;
      RECT 10.83 0.32 11.915 0.51 ;
      RECT 10.83 0.32 11.02 0.945 ;
      RECT 9.14 0.755 11.02 0.945 ;
      RECT 7.125 0.32 7.315 0.97 ;
      RECT 7.035 0.78 7.315 0.97 ;
      RECT 11.725 0.32 11.915 1.21 ;
      RECT 11.725 1.02 14.35 1.21 ;
      RECT 9.14 0.32 9.33 1.335 ;
      RECT 9.05 1.145 9.33 1.335 ;
      RECT 8.105 0.32 8.295 2.16 ;
      RECT 6.935 1.97 8.295 2.16 ;
      RECT 14.16 1.02 14.35 2.375 ;
      RECT 6.935 1.97 7.125 2.65 ;
      RECT 6.845 2.46 7.125 2.65 ;
      RECT 13.77 0.585 14.765 0.775 ;
      RECT 14.575 1.81 15.775 2 ;
      RECT 14.575 0.585 14.765 2.765 ;
      RECT 13.74 2.575 14.765 2.765 ;
      RECT 16.105 0.345 16.295 1.21 ;
      RECT 15.095 1.02 16.295 1.21 ;
      RECT 15.975 1.02 16.165 2.48 ;
  END
END SDQV2_7TV50

MACRO SDRNQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDRNQV1_7TV50 0 0 ;
  SIZE 18.24 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.615 1.56 6.16 1.825 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.95 2.41 2.34 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 17.75 0.445 17.94 2.48 ;
        RECT 17.75 0.445 18.12 0.88 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.665 1.52 9.96 2.15 ;
        RECT 9.665 1.96 12.205 2.15 ;
        RECT 12.015 1.96 12.205 2.925 ;
        RECT 14.54 1.81 14.73 2.925 ;
        RECT 12.015 2.735 14.73 2.925 ;
        RECT 14.54 1.81 15.625 2 ;
    END
  END RDN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.6 1.04 3.41 1.23 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.68 1.36 ;
        RECT 4.08 1.125 4.68 1.36 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.42 1.285 3.48 ;
        RECT 4.265 2.965 4.545 3.48 ;
        RECT 10.055 2.74 10.335 3.48 ;
        RECT 11.555 2.35 11.79 3.48 ;
        RECT 14.97 2.36 15.25 3.48 ;
        RECT 16.79 2.36 17.07 3.48 ;
        RECT 0 3.24 18.24 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.82 ;
        RECT 4.455 -0.12 4.735 0.82 ;
        RECT 5.945 -0.12 6.225 0.82 ;
        RECT 10.965 -0.12 11.245 0.98 ;
        RECT 14.52 -0.12 14.8 0.78 ;
        RECT 16.81 -0.12 17.09 0.74 ;
        RECT 0 -0.12 18.24 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.66 1.46 ;
        RECT -0.12 -0.24 18.36 1.405 ;
        RECT 7.56 -0.24 14.515 1.565 ;
        RECT 7.56 -0.24 18.36 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.66 1.405 7.56 3.94 ;
        RECT -0.58 1.46 7.56 3.94 ;
        RECT 14.515 1.46 18.82 3.94 ;
        RECT -0.58 1.565 18.82 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.56 3.215 1.75 ;
      RECT 3.025 1.56 3.215 2.185 ;
      RECT 0.2 0.54 0.39 2.645 ;
      RECT 5.08 1.02 6.615 1.21 ;
      RECT 5.08 0.54 5.28 2.375 ;
      RECT 5.08 2.185 5.42 2.375 ;
      RECT 6.89 1.42 7.225 1.7 ;
      RECT 6.89 0.54 7.08 2.375 ;
      RECT 6.795 2.185 7.08 2.375 ;
      RECT 2.755 0.585 3.805 0.775 ;
      RECT 2.65 2.42 2.84 2.765 ;
      RECT 3.615 0.585 3.805 2.765 ;
      RECT 7.48 0.54 7.67 2.765 ;
      RECT 2.65 2.575 7.67 2.765 ;
      RECT 9.135 0.745 9.525 0.935 ;
      RECT 9.135 0.745 9.325 2.54 ;
      RECT 9.135 2.35 11.245 2.54 ;
      RECT 8.39 0.355 10.38 0.545 ;
      RECT 10.19 0.355 10.38 1.37 ;
      RECT 10.19 1.18 11.62 1.37 ;
      RECT 8.39 0.355 8.58 2.535 ;
      RECT 8.285 2.345 8.58 2.535 ;
      RECT 11.91 0.7 12.1 1.76 ;
      RECT 10.59 1.57 12.595 1.76 ;
      RECT 12.405 1.57 12.595 2.535 ;
      RECT 12.405 2.345 12.685 2.535 ;
      RECT 12.39 1.18 13.15 1.37 ;
      RECT 12.96 1.18 13.15 2.1 ;
      RECT 12.96 1.91 13.91 2.1 ;
      RECT 12.765 0.745 14.3 0.935 ;
      RECT 14.11 0.98 16.065 1.17 ;
      RECT 14.11 0.745 14.3 2.535 ;
      RECT 13.255 2.345 14.3 2.535 ;
      RECT 16.265 0.5 16.455 1.61 ;
      RECT 14.535 1.42 17.51 1.61 ;
      RECT 15.865 1.42 16.055 2.48 ;
  END
END SDRNQV1_7TV50

MACRO SDRNQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDRNQV2_7TV50 0 0 ;
  SIZE 19.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.615 1.56 6.16 1.825 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.95 2.41 2.34 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 17.75 0.445 17.94 2.48 ;
        RECT 17.75 0.445 18.12 0.88 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.665 1.52 9.96 2.15 ;
        RECT 9.665 1.96 12.205 2.15 ;
        RECT 12.015 1.96 12.205 2.925 ;
        RECT 14.54 1.81 14.73 2.925 ;
        RECT 12.015 2.735 14.73 2.925 ;
        RECT 14.54 1.81 15.525 2 ;
    END
  END RDN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.6 1.04 3.41 1.23 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.68 1.36 ;
        RECT 4.08 1.125 4.68 1.36 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.42 1.285 3.48 ;
        RECT 4.265 2.965 4.545 3.48 ;
        RECT 5.885 2.965 6.165 3.48 ;
        RECT 10.055 2.74 10.335 3.48 ;
        RECT 11.555 2.35 11.79 3.48 ;
        RECT 14.97 2.36 15.25 3.48 ;
        RECT 16.79 2.36 17.07 3.48 ;
        RECT 18.555 2.2 18.835 3.48 ;
        RECT 0 3.24 19.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.82 ;
        RECT 4.455 -0.12 4.735 0.82 ;
        RECT 5.945 -0.12 6.225 0.82 ;
        RECT 10.965 -0.12 11.245 0.98 ;
        RECT 14.52 -0.12 14.8 0.78 ;
        RECT 16.81 -0.12 17.09 0.74 ;
        RECT 18.61 -0.12 18.89 0.725 ;
        RECT 0 -0.12 19.2 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.66 1.46 ;
        RECT -0.12 -0.24 19.32 1.405 ;
        RECT 7.56 -0.24 14.515 1.565 ;
        RECT 7.56 -0.24 19.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.66 1.405 7.56 3.94 ;
        RECT -0.58 1.46 7.56 3.94 ;
        RECT 14.515 1.46 19.78 3.94 ;
        RECT -0.58 1.565 19.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.56 3.215 1.75 ;
      RECT 3.025 1.56 3.215 2.185 ;
      RECT 0.2 0.54 0.39 2.645 ;
      RECT 5.08 1.02 6.615 1.21 ;
      RECT 5.08 0.54 5.28 2.375 ;
      RECT 5.08 2.185 5.42 2.375 ;
      RECT 6.89 1.42 7.225 1.7 ;
      RECT 6.89 0.54 7.08 2.375 ;
      RECT 6.795 2.185 7.08 2.375 ;
      RECT 2.755 0.585 3.805 0.775 ;
      RECT 2.65 2.42 2.84 2.765 ;
      RECT 3.615 0.585 3.805 2.765 ;
      RECT 7.48 0.54 7.67 2.765 ;
      RECT 2.65 2.575 7.67 2.765 ;
      RECT 9.135 0.745 9.525 0.935 ;
      RECT 9.135 0.745 9.325 2.54 ;
      RECT 9.135 2.35 11.245 2.54 ;
      RECT 8.39 0.355 10.38 0.545 ;
      RECT 10.19 0.355 10.38 1.37 ;
      RECT 10.19 1.18 11.62 1.37 ;
      RECT 8.39 0.355 8.58 2.535 ;
      RECT 8.285 2.345 8.58 2.535 ;
      RECT 11.91 0.7 12.1 1.76 ;
      RECT 10.59 1.57 12.595 1.76 ;
      RECT 12.405 1.57 12.595 2.535 ;
      RECT 12.405 2.345 12.685 2.535 ;
      RECT 12.39 1.18 13.15 1.37 ;
      RECT 12.96 1.18 13.15 2.1 ;
      RECT 12.96 1.91 13.91 2.1 ;
      RECT 12.765 0.745 14.3 0.935 ;
      RECT 14.11 0.98 16.065 1.17 ;
      RECT 14.11 0.745 14.3 2.535 ;
      RECT 13.255 2.345 14.3 2.535 ;
      RECT 16.265 1.075 17.465 1.265 ;
      RECT 16.265 0.5 16.455 1.61 ;
      RECT 14.535 1.42 16.455 1.61 ;
      RECT 15.865 1.42 16.055 2.48 ;
  END
END SDRNQV2_7TV50

MACRO SDRQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDRQV1_7TV50 0 0 ;
  SIZE 19.2 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.76 1.56 6.36 1.8 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.945 2.41 2.335 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 18.475 0.56 18.665 2.48 ;
        RECT 18.475 0.56 19.08 0.88 ;
    END
  END Q
  PIN RD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.52 2.48 14.76 3 ;
        RECT 14.52 2.81 14.9 3 ;
    END
  END RD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.265 ;
        RECT 0.6 1.075 3.41 1.265 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.08 1.605 4.68 1.84 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.51 1.285 3.48 ;
        RECT 4.265 2.925 4.5 3.48 ;
        RECT 9.885 2.335 10.165 3.48 ;
        RECT 15.14 2.33 15.375 3.48 ;
        RECT 17.58 2.28 17.86 3.48 ;
        RECT 0 3.24 19.2 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.835 ;
        RECT 4.455 -0.12 4.69 0.795 ;
        RECT 10.285 -0.12 10.565 0.51 ;
        RECT 15.37 -0.12 15.65 0.74 ;
        RECT 17.76 -0.12 18.04 0.58 ;
        RECT 0 -0.12 19.2 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.83 -0.24 7.72 1.6 ;
        RECT 9.925 -0.24 14.145 1.545 ;
        RECT 12.525 -0.24 14.145 1.565 ;
        RECT -0.12 -0.24 19.32 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.83 3.94 ;
        RECT 7.72 1.46 9.925 3.94 ;
        RECT 7.72 1.545 12.525 3.94 ;
        RECT 7.72 1.565 19.78 3.94 ;
        RECT 14.145 1.46 19.78 3.94 ;
        RECT -0.58 1.6 19.78 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.485 3.215 1.675 ;
      RECT 3.025 1.485 3.215 2.18 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.28 2.025 6.65 2.215 ;
      RECT 5.28 0.735 5.47 2.65 ;
      RECT 5.19 2.46 5.47 2.65 ;
      RECT 7.035 0.78 7.315 0.97 ;
      RECT 7.035 0.78 7.225 2.65 ;
      RECT 6.845 2.46 7.225 2.65 ;
      RECT 2.65 2.355 2.84 2.72 ;
      RECT 2.65 2.53 4.89 2.72 ;
      RECT 4.7 2.53 4.89 3.04 ;
      RECT 7.48 2.615 7.67 3.04 ;
      RECT 4.7 2.85 7.67 3.04 ;
      RECT 4.89 0.345 7.86 0.535 ;
      RECT 7.67 0.345 7.86 0.745 ;
      RECT 2.755 0.56 3.875 0.75 ;
      RECT 3.685 0.56 3.875 1.185 ;
      RECT 4.89 0.345 5.08 1.185 ;
      RECT 3.685 0.995 5.08 1.185 ;
      RECT 8.57 1.52 11.39 1.71 ;
      RECT 8.57 0.54 8.76 2.57 ;
      RECT 8.285 2.38 8.76 2.57 ;
      RECT 7.895 1.02 8.28 1.21 ;
      RECT 9.145 1.91 12.14 2.1 ;
      RECT 7.895 1.02 8.085 3.005 ;
      RECT 9.145 1.91 9.335 3.005 ;
      RECT 7.895 2.815 9.335 3.005 ;
      RECT 12.71 0.745 12.99 0.935 ;
      RECT 11.245 0.725 11.525 1.32 ;
      RECT 12.71 0.745 12.9 1.32 ;
      RECT 9.85 1.13 12.9 1.32 ;
      RECT 12.34 1.13 12.53 2.565 ;
      RECT 11.485 2.375 12.53 2.565 ;
      RECT 10.83 0.32 13.38 0.51 ;
      RECT 10.83 0.32 11.02 0.93 ;
      RECT 9.095 0.74 11.02 0.93 ;
      RECT 9.095 0.74 9.285 1.255 ;
      RECT 13.19 0.32 13.38 1.415 ;
      RECT 13.58 0.545 13.95 0.735 ;
      RECT 16.315 0.5 16.505 1.36 ;
      RECT 13.58 1.17 17.515 1.36 ;
      RECT 13.58 0.545 13.77 2.52 ;
      RECT 12.73 2.33 13.77 2.52 ;
      RECT 12.73 2.33 12.92 2.61 ;
      RECT 16.905 0.415 17.095 0.97 ;
      RECT 16.905 0.78 17.905 0.97 ;
      RECT 17.715 0.78 17.905 1.93 ;
      RECT 13.97 1.74 18.235 1.93 ;
      RECT 16.775 1.74 16.965 2.48 ;
  END
END SDRQV1_7TV50

MACRO SDRQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDRQV2_7TV50 0 0 ;
  SIZE 20.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.76 1.56 6.36 1.8 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.945 2.41 2.335 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 18.475 0.56 18.665 2.48 ;
        RECT 18.475 0.56 19.08 0.88 ;
    END
  END Q
  PIN RD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 14.52 2.48 14.76 3 ;
        RECT 14.52 2.81 14.9 3 ;
    END
  END RD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 0.56 0.84 1.265 ;
        RECT 0.6 1.075 3.41 1.265 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.52 4.68 1.84 ;
        RECT 4.08 1.605 4.68 1.84 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.51 1.285 3.48 ;
        RECT 4.265 2.925 4.5 3.48 ;
        RECT 9.885 2.335 10.165 3.48 ;
        RECT 15.14 2.33 15.375 3.48 ;
        RECT 17.58 2.28 17.86 3.48 ;
        RECT 19.28 2.28 19.56 3.48 ;
        RECT 0 3.24 20.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.835 ;
        RECT 4.455 -0.12 4.69 0.795 ;
        RECT 6.135 -0.12 6.415 0.97 ;
        RECT 10.285 -0.12 10.565 0.51 ;
        RECT 15.37 -0.12 15.65 0.74 ;
        RECT 17.76 -0.12 18.04 0.58 ;
        RECT 19.56 -0.12 19.84 0.725 ;
        RECT 0 -0.12 20.16 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.83 -0.24 7.72 1.6 ;
        RECT 9.925 -0.24 14.145 1.545 ;
        RECT 12.525 -0.24 14.145 1.565 ;
        RECT -0.12 -0.24 20.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.83 3.94 ;
        RECT 7.72 1.46 9.925 3.94 ;
        RECT 7.72 1.545 12.525 3.94 ;
        RECT 7.72 1.565 20.74 3.94 ;
        RECT 14.145 1.46 20.74 3.94 ;
        RECT -0.58 1.6 20.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.485 3.215 1.675 ;
      RECT 3.025 1.485 3.215 2.18 ;
      RECT 0.2 0.595 0.39 2.475 ;
      RECT 5.28 2.025 6.65 2.215 ;
      RECT 5.28 0.735 5.47 2.65 ;
      RECT 5.19 2.46 5.47 2.65 ;
      RECT 7.035 0.78 7.315 0.97 ;
      RECT 7.035 0.78 7.225 2.65 ;
      RECT 6.845 2.46 7.225 2.65 ;
      RECT 2.65 2.355 2.84 2.72 ;
      RECT 2.65 2.53 4.89 2.72 ;
      RECT 4.7 2.53 4.89 3.04 ;
      RECT 7.48 2.615 7.67 3.04 ;
      RECT 4.7 2.85 7.67 3.04 ;
      RECT 4.89 0.345 5.935 0.535 ;
      RECT 6.615 0.39 7.86 0.58 ;
      RECT 7.67 0.39 7.86 0.745 ;
      RECT 2.755 0.56 3.875 0.75 ;
      RECT 3.685 0.56 3.875 1.185 ;
      RECT 5.745 0.345 5.935 1.36 ;
      RECT 4.89 0.345 5.08 1.185 ;
      RECT 3.685 0.995 5.08 1.185 ;
      RECT 6.615 0.39 6.805 1.36 ;
      RECT 5.745 1.17 6.805 1.36 ;
      RECT 8.57 1.52 11.39 1.71 ;
      RECT 8.57 0.54 8.76 2.57 ;
      RECT 8.285 2.38 8.76 2.57 ;
      RECT 7.895 1.02 8.28 1.21 ;
      RECT 9.145 1.91 12.14 2.1 ;
      RECT 7.895 1.02 8.085 3.005 ;
      RECT 9.145 1.91 9.335 3.005 ;
      RECT 7.895 2.815 9.335 3.005 ;
      RECT 12.71 0.745 12.99 0.935 ;
      RECT 11.245 0.725 11.525 1.32 ;
      RECT 12.71 0.745 12.9 1.32 ;
      RECT 9.85 1.13 12.9 1.32 ;
      RECT 12.34 1.13 12.53 2.565 ;
      RECT 11.485 2.375 12.53 2.565 ;
      RECT 10.83 0.32 13.38 0.51 ;
      RECT 10.83 0.32 11.02 0.93 ;
      RECT 9.095 0.74 11.02 0.93 ;
      RECT 9.095 0.74 9.285 1.255 ;
      RECT 13.19 0.32 13.38 1.415 ;
      RECT 13.58 0.545 13.95 0.735 ;
      RECT 16.315 0.5 16.505 1.36 ;
      RECT 13.58 1.17 17.515 1.36 ;
      RECT 13.58 0.545 13.77 2.52 ;
      RECT 12.73 2.33 13.77 2.52 ;
      RECT 12.73 2.33 12.92 2.61 ;
      RECT 16.905 0.415 17.095 0.97 ;
      RECT 16.905 0.78 17.905 0.97 ;
      RECT 17.715 0.78 17.905 1.93 ;
      RECT 13.97 1.74 18.235 1.93 ;
      RECT 16.775 1.74 16.965 2.48 ;
  END
END SDRQV2_7TV50

MACRO SDSRNQV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDSRNQV1_7TV50 0 0 ;
  SIZE 20.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.56 1.08 6.16 1.32 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.95 2.41 2.34 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 19.28 0.6 19.895 0.84 ;
        RECT 19.705 0.6 19.895 2.48 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.475 2.31 11.665 2.775 ;
        RECT 9.185 2.585 11.665 2.775 ;
        RECT 11.475 2.31 12.555 2.5 ;
        RECT 12.365 2.31 12.555 2.985 ;
        RECT 18.36 1.845 18.6 2.985 ;
        RECT 12.365 2.795 18.6 2.985 ;
    END
  END RDN
  PIN SDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.03 0.32 12.22 1.1 ;
        RECT 11.94 0.91 12.22 1.1 ;
        RECT 12.03 0.32 15.48 0.51 ;
        RECT 15.29 0.32 15.48 1.36 ;
        RECT 15.29 1.04 15.72 1.36 ;
    END
  END SDN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.6 1.04 3.41 1.23 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.68 1.36 ;
        RECT 4.08 1.125 4.68 1.36 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.38 1.285 3.48 ;
        RECT 4.265 2.965 4.545 3.48 ;
        RECT 11.865 2.7 12.145 3.48 ;
        RECT 18.81 2.28 19.09 3.48 ;
        RECT 0 3.24 20.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.81 ;
        RECT 4.455 -0.12 4.735 0.82 ;
        RECT 5.945 -0.12 6.225 0.765 ;
        RECT 10.845 -0.12 11.125 0.7 ;
        RECT 16.42 -0.12 16.7 0.875 ;
        RECT 18.71 -0.12 18.99 0.83 ;
        RECT 0 -0.12 20.16 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.66 1.46 ;
        RECT -0.12 -0.24 5.015 1.405 ;
        RECT -0.12 -0.24 20.28 1.35 ;
        RECT 12.52 -0.24 15.245 1.565 ;
        RECT 12.52 -0.24 20.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.66 1.405 12.52 3.94 ;
        RECT 5.015 1.35 12.52 3.94 ;
        RECT -0.58 1.46 12.52 3.94 ;
        RECT 15.245 1.46 20.74 3.94 ;
        RECT -0.58 1.565 20.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.56 3.215 1.75 ;
      RECT 3.025 1.56 3.215 2.185 ;
      RECT 0.2 0.54 0.39 2.62 ;
      RECT 5.09 1.75 6.16 1.94 ;
      RECT 5.09 0.485 5.29 2.375 ;
      RECT 5.01 2.185 5.29 2.375 ;
      RECT 6.585 0.53 7.125 0.72 ;
      RECT 6.585 0.53 6.775 2.375 ;
      RECT 6.345 2.185 6.775 2.375 ;
      RECT 2.755 0.585 3.805 0.775 ;
      RECT 7.48 0.43 7.67 1.375 ;
      RECT 7.045 1.185 7.67 1.375 ;
      RECT 2.65 2.34 2.84 2.765 ;
      RECT 3.615 0.585 3.805 2.765 ;
      RECT 7.045 1.185 7.235 2.765 ;
      RECT 2.65 2.575 7.235 2.765 ;
      RECT 8.7 2.135 10.645 2.325 ;
      RECT 8.39 0.43 8.58 1.105 ;
      RECT 7.895 0.915 11.5 1.105 ;
      RECT 7.895 0.915 8.085 2.365 ;
      RECT 12.555 1.215 12.745 1.495 ;
      RECT 8.87 1.305 12.745 1.495 ;
      RECT 12.945 0.71 13.245 0.9 ;
      RECT 10.12 1.695 13.135 1.885 ;
      RECT 11.045 1.695 11.235 2.32 ;
      RECT 10.955 2.13 11.235 2.32 ;
      RECT 12.945 0.71 13.135 2.595 ;
      RECT 12.775 2.405 13.135 2.595 ;
      RECT 13.335 1.145 14.52 1.335 ;
      RECT 13.335 1.145 13.525 2.205 ;
      RECT 16.29 2.3 16.48 2.595 ;
      RECT 14.475 2.405 16.48 2.595 ;
      RECT 13.865 0.71 14.91 0.9 ;
      RECT 14.72 0.71 14.91 2 ;
      RECT 13.725 1.81 17.705 2 ;
      RECT 13.725 1.81 13.915 2.595 ;
      RECT 13.625 2.405 13.915 2.595 ;
      RECT 17.055 0.595 17.245 1.265 ;
      RECT 16.42 1.075 19.365 1.265 ;
      RECT 17.945 1.075 18.135 2.56 ;
  END
END SDSRNQV1_7TV50

MACRO SDSRNQV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDSRNQV2_7TV50 0 0 ;
  SIZE 21.12 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 5.56 1.08 6.16 1.32 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.04 1.95 2.41 2.34 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 19.28 0.6 19.895 0.84 ;
        RECT 19.705 0.6 19.895 2.48 ;
    END
  END Q
  PIN RDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.475 2.31 11.665 2.775 ;
        RECT 9.185 2.585 11.665 2.775 ;
        RECT 11.475 2.31 12.555 2.5 ;
        RECT 12.365 2.31 12.555 2.985 ;
        RECT 18.36 1.845 18.6 2.985 ;
        RECT 12.365 2.795 18.6 2.985 ;
    END
  END RDN
  PIN SDN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.03 0.32 12.22 1.1 ;
        RECT 11.94 0.91 12.22 1.1 ;
        RECT 12.03 0.32 15.48 0.51 ;
        RECT 15.29 0.32 15.48 1.36 ;
        RECT 15.29 1.04 15.72 1.36 ;
    END
  END SDN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.04 0.84 1.36 ;
        RECT 0.6 1.04 3.41 1.23 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.44 1.04 4.68 1.36 ;
        RECT 4.08 1.125 4.68 1.36 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.005 2.38 1.285 3.48 ;
        RECT 4.265 2.965 4.545 3.48 ;
        RECT 11.865 2.7 12.145 3.48 ;
        RECT 18.81 2.28 19.09 3.48 ;
        RECT 20.51 2.28 20.79 3.48 ;
        RECT 0 3.24 21.12 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.81 ;
        RECT 4.455 -0.12 4.735 0.82 ;
        RECT 5.945 -0.12 6.225 0.765 ;
        RECT 10.845 -0.12 11.125 0.7 ;
        RECT 16.42 -0.12 16.7 0.875 ;
        RECT 18.71 -0.12 18.99 0.83 ;
        RECT 20.51 -0.12 20.79 0.75 ;
        RECT 0 -0.12 21.12 0.12 ;
    END
  END VSS
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT -0.12 -0.24 2.66 1.46 ;
        RECT -0.12 -0.24 5.015 1.405 ;
        RECT -0.12 -0.24 21.24 1.35 ;
        RECT 12.52 -0.24 15.245 1.565 ;
        RECT 12.52 -0.24 21.24 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT 2.66 1.405 12.52 3.94 ;
        RECT 5.015 1.35 12.52 3.94 ;
        RECT -0.58 1.46 12.52 3.94 ;
        RECT 15.245 1.46 21.7 3.94 ;
        RECT -0.58 1.565 21.7 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.56 3.215 1.75 ;
      RECT 3.025 1.56 3.215 2.185 ;
      RECT 0.2 0.54 0.39 2.62 ;
      RECT 5.09 1.75 6.16 1.94 ;
      RECT 5.09 0.485 5.29 2.375 ;
      RECT 5.01 2.185 5.29 2.375 ;
      RECT 6.585 0.53 7.125 0.72 ;
      RECT 6.585 0.53 6.775 2.375 ;
      RECT 6.345 2.185 6.775 2.375 ;
      RECT 2.755 0.585 3.805 0.775 ;
      RECT 7.48 0.43 7.67 1.33 ;
      RECT 7.045 1.14 7.67 1.33 ;
      RECT 2.65 2.34 2.84 2.765 ;
      RECT 3.615 0.585 3.805 2.765 ;
      RECT 7.045 1.14 7.235 2.765 ;
      RECT 2.65 2.575 7.235 2.765 ;
      RECT 8.7 2.135 10.645 2.325 ;
      RECT 8.39 0.43 8.58 1.105 ;
      RECT 7.895 0.915 11.5 1.105 ;
      RECT 7.895 0.915 8.085 2.365 ;
      RECT 12.555 1.215 12.745 1.495 ;
      RECT 8.87 1.305 12.745 1.495 ;
      RECT 12.945 0.71 13.245 0.9 ;
      RECT 10.12 1.695 13.135 1.885 ;
      RECT 11 1.695 11.19 2.32 ;
      RECT 10.955 2.13 11.235 2.32 ;
      RECT 12.945 0.71 13.135 2.595 ;
      RECT 12.775 2.405 13.135 2.595 ;
      RECT 13.335 1.145 14.52 1.335 ;
      RECT 13.335 1.145 13.525 2.205 ;
      RECT 16.29 2.3 16.48 2.595 ;
      RECT 14.475 2.405 16.48 2.595 ;
      RECT 13.865 0.71 14.91 0.9 ;
      RECT 14.72 0.71 14.91 2 ;
      RECT 13.725 1.81 17.705 2 ;
      RECT 13.725 1.81 13.915 2.595 ;
      RECT 13.625 2.405 13.915 2.595 ;
      RECT 17.055 0.595 17.245 1.265 ;
      RECT 16.42 1.075 19.365 1.265 ;
      RECT 17.945 1.075 18.135 2.56 ;
  END
END SDSRNQV2_7TV50

MACRO TBUFV1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFV1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 1.88 0.975 2.28 ;
    END
  END I
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 1.04 2.995 1.38 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.155 2.97 1.435 3.48 ;
        RECT 5.435 2.7 5.715 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.155 -0.12 1.435 0.39 ;
        RECT 5.045 -0.12 5.325 0.675 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.24 0.39 6.6 0.58 ;
        RECT 6.36 1.52 6.6 1.84 ;
        RECT 6.41 0.39 6.6 2.5 ;
        RECT 6.285 2.31 6.6 2.5 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.915 -0.24 4.97 1.53 ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.915 3.94 ;
        RECT 4.97 1.46 7.3 3.94 ;
        RECT -0.58 1.53 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.245 2.56 0.525 2.77 ;
      RECT 0.245 2.58 2.84 2.77 ;
      RECT 2.56 2.58 2.84 3.025 ;
      RECT 4.085 0.71 4.43 0.9 ;
      RECT 1.845 0.98 2.035 1.99 ;
      RECT 1.845 1.8 4.43 1.99 ;
      RECT 4.24 0.71 4.43 2.545 ;
      RECT 0.195 0.59 2.455 0.78 ;
      RECT 5.045 1.515 5.52 1.705 ;
      RECT 1.38 0.59 1.57 2.38 ;
      RECT 1.38 2.19 3.84 2.38 ;
      RECT 3.65 2.19 3.84 2.935 ;
      RECT 5.045 1.515 5.235 2.935 ;
      RECT 3.65 2.745 5.235 2.935 ;
      RECT 3.205 0.32 4.845 0.51 ;
      RECT 3.205 0.32 3.395 0.825 ;
      RECT 4.655 0.32 4.845 1.29 ;
      RECT 4.655 1.1 6.045 1.29 ;
      RECT 5.855 1.1 6.045 2.04 ;
  END
END TBUFV1_7TV50

MACRO TBUFV2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFV2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.49 1.91 0.92 2.32 ;
    END
  END I
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.52 1.04 2.98 1.36 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.125 2.925 1.405 3.48 ;
        RECT 5.735 2.31 6.015 3.48 ;
        RECT 7.435 2.385 7.715 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.17 -0.12 1.36 0.435 ;
        RECT 5.06 -0.12 5.25 0.66 ;
        RECT 7.485 -0.12 7.675 0.66 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.54 0.425 6.82 0.615 ;
        RECT 6.63 0.425 6.82 2.545 ;
        RECT 6.63 1.56 7.12 1.8 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.7 -0.24 4.895 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.7 3.94 ;
        RECT 4.895 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.215 2.535 2.265 2.725 ;
      RECT 2.075 2.535 2.265 3.04 ;
      RECT 2.075 2.85 3.8 3.04 ;
      RECT 1.63 1.06 1.82 1.82 ;
      RECT 4.055 0.71 4.335 1.82 ;
      RECT 1.63 1.63 4.58 1.82 ;
      RECT 4.39 1.63 4.58 2.545 ;
      RECT 0.21 0.58 0.4 0.86 ;
      RECT 2.13 0.58 2.32 0.86 ;
      RECT 0.21 0.66 2.32 0.86 ;
      RECT 5.24 1.35 5.67 1.54 ;
      RECT 1.24 0.66 1.43 2.335 ;
      RECT 1.24 2.145 2.655 2.335 ;
      RECT 2.465 2.145 2.655 2.535 ;
      RECT 2.465 2.345 4.19 2.535 ;
      RECT 4 2.345 4.19 2.935 ;
      RECT 5.24 1.35 5.43 2.935 ;
      RECT 4 2.745 5.43 2.935 ;
      RECT 3.09 0.32 4.86 0.51 ;
      RECT 3.09 0.32 3.28 0.86 ;
      RECT 4.67 0.32 4.86 1.1 ;
      RECT 4.67 0.91 6.385 1.1 ;
      RECT 6.195 0.91 6.385 2.045 ;
  END
END TBUFV2_7TV50

MACRO TBUFV3_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFV3_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.49 1.48 0.89 1.84 ;
    END
  END I
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.39 1.035 2.8 1.395 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.195 2.97 1.475 3.48 ;
        RECT 5.145 2.39 5.425 3.48 ;
        RECT 6.845 2.355 7.125 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.83 ;
        RECT 4.665 -0.12 4.945 0.39 ;
        RECT 6.525 -0.12 6.805 0.615 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.67 0.56 6.23 0.84 ;
        RECT 6.04 0.56 6.23 2.545 ;
        RECT 7.47 0.56 7.66 1.8 ;
        RECT 6.04 1.56 7.96 1.8 ;
        RECT 7.77 1.56 7.96 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.47 -0.24 4.375 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.47 3.94 ;
        RECT 4.375 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.205 2.58 2.155 2.77 ;
      RECT 1.965 2.76 3.74 2.955 ;
      RECT 3.55 2.76 3.74 3.04 ;
      RECT 1.48 1.42 1.76 1.61 ;
      RECT 1.57 1.42 1.76 1.99 ;
      RECT 3.645 0.71 3.925 1.99 ;
      RECT 1.57 1.8 4.53 1.99 ;
      RECT 4.34 1.8 4.53 2.545 ;
      RECT 0.2 0.595 0.39 1.22 ;
      RECT 2 0.595 2.19 1.22 ;
      RECT 0.2 1.03 2.19 1.22 ;
      RECT 4.755 1.04 5.08 1.23 ;
      RECT 1.09 1.03 1.28 2.38 ;
      RECT 1.09 2.19 2.545 2.38 ;
      RECT 2.355 2.37 4.13 2.56 ;
      RECT 3.94 2.37 4.13 3.015 ;
      RECT 4.755 1.04 4.945 3.015 ;
      RECT 3.94 2.825 4.945 3.015 ;
      RECT 2.855 0.32 4.315 0.51 ;
      RECT 4.125 0.32 4.315 0.825 ;
      RECT 4.125 0.635 5.47 0.825 ;
      RECT 2.855 0.32 3.135 0.83 ;
      RECT 5.28 0.635 5.47 1.995 ;
      RECT 5.28 1.805 5.815 1.995 ;
  END
END TBUFV3_7TV50

MACRO TBUFV4_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFV4_7TV50 0 0 ;
  SIZE 10.08 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.73 1.585 1.36 1.775 ;
        RECT 1.04 1.56 1.36 1.8 ;
        RECT 1.04 1.575 1.815 1.765 ;
    END
  END I
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.84 1.08 4.3 1.395 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.255 2.65 0.535 3.48 ;
        RECT 2.015 2.97 2.295 3.48 ;
        RECT 6.165 2.325 6.445 3.48 ;
        RECT 7.895 2.405 8.175 3.48 ;
        RECT 9.595 2.405 9.875 3.48 ;
        RECT 0 3.24 10.08 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.735 ;
        RECT 1.955 -0.12 2.235 0.82 ;
        RECT 5.64 -0.12 5.92 0.39 ;
        RECT 7.5 -0.12 7.78 0.65 ;
        RECT 9.3 -0.12 9.58 0.65 ;
        RECT 0 -0.12 10.08 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.645 0.595 7.25 0.875 ;
        RECT 7.06 0.595 7.25 2.475 ;
        RECT 7.06 1.08 7.6 1.32 ;
        RECT 8.445 0.595 8.635 1.27 ;
        RECT 7.06 1.08 8.98 1.27 ;
        RECT 8.79 1.08 8.98 2.475 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 3.76 -0.24 5.535 1.53 ;
        RECT -0.12 -0.24 10.2 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 3.76 3.94 ;
        RECT 5.535 1.46 10.66 3.94 ;
        RECT -0.58 1.53 10.66 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.105 2.58 3.035 2.77 ;
      RECT 2.845 2.58 3.035 2.98 ;
      RECT 2.845 2.79 4.71 2.98 ;
      RECT 4.43 2.79 4.71 3.04 ;
      RECT 2.525 1.41 2.715 1.99 ;
      RECT 4.62 0.71 4.9 1.99 ;
      RECT 2.525 1.8 5.49 1.99 ;
      RECT 5.3 1.8 5.49 2.545 ;
      RECT 1.1 0.585 1.29 1.21 ;
      RECT 2.9 0.585 3.09 1.21 ;
      RECT 1.1 1.02 3.09 1.21 ;
      RECT 5.775 1.03 6.055 1.31 ;
      RECT 2.12 1.02 2.31 2.38 ;
      RECT 2.12 2.19 4.03 2.38 ;
      RECT 3.84 2.34 5.1 2.53 ;
      RECT 4.91 2.34 5.1 2.935 ;
      RECT 5.775 1.03 5.965 2.935 ;
      RECT 4.91 2.745 5.965 2.935 ;
      RECT 3.86 0.32 5.375 0.51 ;
      RECT 5.185 0.32 5.375 0.78 ;
      RECT 5.185 0.59 6.445 0.78 ;
      RECT 3.86 0.32 4.05 0.865 ;
      RECT 6.255 0.59 6.445 1.995 ;
      RECT 6.255 1.805 6.835 1.995 ;
  END
END TBUFV4_7TV50

MACRO XNOR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2V1_7TV50 0 0 ;
  SIZE 5.28 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.455 1.1 2.8 1.29 ;
        RECT 2.545 1.08 2.735 1.915 ;
        RECT 2.48 1.08 2.8 1.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.44 1.06 4.06 1.32 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.235 2.405 0.515 3.48 ;
        RECT 3.905 2.745 4.185 3.48 ;
        RECT 0 3.24 5.28 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.235 -0.12 0.475 0.61 ;
        RECT 3.855 -0.12 4.135 0.565 ;
        RECT 0 -0.12 5.28 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.065 0.71 1.255 2.73 ;
        RECT 1.52 2.52 1.84 2.76 ;
        RECT 1.065 2.54 2.115 2.73 ;
        RECT 1.065 0.71 2.275 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.62 -0.24 2.59 1.545 ;
        RECT -0.12 -0.24 5.4 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.62 3.94 ;
        RECT 2.59 1.46 5.86 3.94 ;
        RECT -0.58 1.545 5.86 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.675 0.32 3.19 0.51 ;
      RECT 0.675 0.32 0.865 1.295 ;
      RECT 3 0.32 3.19 2.515 ;
      RECT 2.975 2.325 3.255 2.515 ;
      RECT 1.505 1.845 1.695 2.32 ;
      RECT 1.505 2.13 2.595 2.32 ;
      RECT 4.8 0.58 4.99 2.49 ;
      RECT 3.495 2.3 4.99 2.49 ;
      RECT 2.405 2.13 2.595 2.905 ;
      RECT 3.495 2.3 3.685 2.905 ;
      RECT 2.405 2.715 3.685 2.905 ;
  END
END XNOR2V1_7TV50

MACRO XNOR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2V2_7TV50 0 0 ;
  SIZE 7.68 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.41 0.32 3.6 1.38 ;
        RECT 3.41 0.32 4.495 0.51 ;
        RECT 4.305 0.32 4.495 2.08 ;
        RECT 4.305 1.89 4.72 2.08 ;
        RECT 5.895 1.56 6.64 1.805 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.04 1.56 1.36 2 ;
        RECT 0.63 1.81 1.76 2 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.405 0.435 3.48 ;
        RECT 1.955 2.795 2.235 3.48 ;
        RECT 6.325 2.795 6.605 3.48 ;
        RECT 0 3.24 7.68 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.565 ;
        RECT 1.955 -0.12 2.235 0.565 ;
        RECT 6.275 -0.12 6.555 0.565 ;
        RECT 0 -0.12 7.68 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.48 2 4.05 2.32 ;
        RECT 3.855 0.71 4.05 2.56 ;
        RECT 3.815 0.71 4.095 0.9 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.595 -0.24 5.3 1.53 ;
        RECT -0.12 -0.24 7.8 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.49 3.94 ;
        RECT 5.195 1.46 8.26 3.94 ;
        RECT -0.58 1.53 8.26 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.96 0.665 3.15 2.595 ;
      RECT 1.1 0.525 1.29 0.955 ;
      RECT 1.1 0.765 2.625 0.955 ;
      RECT 4.76 0.455 4.95 1.645 ;
      RECT 1.105 2.36 2.625 2.55 ;
      RECT 2.435 0.765 2.625 2.985 ;
      RECT 4.92 1.455 5.11 2.985 ;
      RECT 2.435 2.795 5.11 2.985 ;
      RECT 5.375 0.375 5.655 0.565 ;
      RECT 5.18 1 5.655 1.205 ;
      RECT 5.465 1.11 7.41 1.3 ;
      RECT 7.22 0.525 7.41 2.48 ;
      RECT 5.465 0.375 5.655 3.03 ;
  END
END XNOR2V2_7TV50

MACRO XNOR3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3V1_7TV50 0 0 ;
  SIZE 11.04 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.545 1.785 1.9 2.38 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.92 0.94 2.365 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.12 1.43 9.52 1.8 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.745 1.345 3.48 ;
        RECT 5.015 2.745 5.295 3.48 ;
        RECT 9.755 2.795 10.035 3.48 ;
        RECT 0 3.24 11.04 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 -0.12 1.345 0.615 ;
        RECT 5.025 -0.12 5.285 0.685 ;
        RECT 9.705 -0.12 9.985 0.615 ;
        RECT 0 -0.12 11.04 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.65 0.56 10.84 2.48 ;
        RECT 10.65 0.56 10.92 0.88 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.74 -0.24 3.81 1.565 ;
        RECT 0.74 -0.24 8.315 1.555 ;
        RECT -0.12 -0.24 11.16 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.74 3.94 ;
        RECT 3.81 1.555 11.62 3.94 ;
        RECT 8.315 1.46 11.62 3.94 ;
        RECT -0.58 1.565 11.62 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.21 1.395 2.455 1.585 ;
      RECT 2.265 1.395 2.455 1.675 ;
      RECT 0.21 0.38 0.4 2.775 ;
      RECT 0.21 2.585 0.495 2.775 ;
      RECT 2.085 0.745 2.845 0.935 ;
      RECT 2.655 1.36 3.84 1.55 ;
      RECT 2.655 0.745 2.845 2.185 ;
      RECT 2.25 1.995 2.845 2.185 ;
      RECT 2.25 1.995 2.44 2.82 ;
      RECT 4.065 0.735 4.345 0.925 ;
      RECT 4.115 0.735 4.345 2.65 ;
      RECT 3.965 2.46 4.345 2.65 ;
      RECT 5.905 0.735 6.265 0.925 ;
      RECT 5.905 0.735 6.105 2.82 ;
      RECT 3.15 0.345 4.81 0.535 ;
      RECT 5.485 0.345 8.21 0.535 ;
      RECT 3.15 0.345 3.34 0.69 ;
      RECT 5.485 0.345 5.675 1.12 ;
      RECT 4.62 0.93 5.675 1.12 ;
      RECT 8.02 0.345 8.21 2.615 ;
      RECT 7.63 2.425 8.21 2.615 ;
      RECT 3.1 2.7 3.29 3.04 ;
      RECT 4.62 0.345 4.81 3.04 ;
      RECT 3.1 2.85 4.81 3.04 ;
      RECT 8.655 0.425 8.945 0.615 ;
      RECT 8.655 0.425 8.845 2.65 ;
      RECT 6.765 0.735 7.285 0.925 ;
      RECT 10.19 1.73 10.38 2.215 ;
      RECT 9.045 2.025 10.38 2.215 ;
      RECT 6.765 0.735 6.955 3.04 ;
      RECT 9.045 2.025 9.235 3.04 ;
      RECT 6.765 2.85 9.235 3.04 ;
  END
END XNOR3V1_7TV50

MACRO XNOR3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3V2_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 0.56 1.8 1.21 ;
        RECT 1.44 0.985 1.8 1.21 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.895 0.95 2.365 ;
        RECT 3.865 1.13 4.055 2.095 ;
        RECT 0.6 1.895 4.055 2.095 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.87 1.26 7.06 2.145 ;
        RECT 7.81 1.1 8 1.45 ;
        RECT 6.87 1.26 8 1.45 ;
        RECT 9.665 1.285 10 1.8 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.765 1.345 3.48 ;
        RECT 5.595 2.745 5.875 3.48 ;
        RECT 10.21 2.795 10.49 3.48 ;
        RECT 12.045 2.405 12.325 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.17 -0.12 1.36 0.66 ;
        RECT 5.65 -0.12 5.84 0.66 ;
        RECT 10.215 -0.12 10.495 0.615 ;
        RECT 12.045 -0.12 12.325 0.615 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.155 0.53 11.4 0.88 ;
        RECT 11.205 0.53 11.4 2.65 ;
    END
  END ZN
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.12 -0.24 9.115 1.555 ;
        RECT -0.12 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.12 3.94 ;
        RECT 9.115 1.46 13.06 3.94 ;
        RECT -0.58 1.555 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.21 0.585 0.505 0.775 ;
      RECT 2.235 1.255 2.8 1.445 ;
      RECT 2.235 1.255 2.425 1.695 ;
      RECT 0.21 1.505 2.425 1.695 ;
      RECT 0.21 0.585 0.4 2.775 ;
      RECT 0.21 2.585 0.49 2.775 ;
      RECT 2.13 0.54 2.32 1.055 ;
      RECT 3.475 0.74 4.445 0.93 ;
      RECT 2.13 0.865 3.665 1.055 ;
      RECT 4.255 0.74 4.445 2.545 ;
      RECT 2.25 2.355 4.445 2.545 ;
      RECT 2.25 2.355 2.44 2.82 ;
      RECT 4.645 0.71 4.925 0.9 ;
      RECT 4.735 0.71 4.925 2.65 ;
      RECT 4.695 2.46 4.975 2.65 ;
      RECT 6.48 0.71 6.845 0.9 ;
      RECT 6.48 0.71 6.67 2.775 ;
      RECT 6.445 2.585 6.725 2.775 ;
      RECT 3.09 0.32 5.39 0.51 ;
      RECT 6.04 0.32 8.79 0.51 ;
      RECT 3.09 0.32 3.28 0.665 ;
      RECT 5.2 1.385 6.23 1.58 ;
      RECT 6.04 0.32 6.23 2.145 ;
      RECT 8.6 0.32 8.79 2.535 ;
      RECT 8.21 2.345 8.79 2.535 ;
      RECT 3.055 2.745 3.335 3.04 ;
      RECT 5.2 0.32 5.39 3.04 ;
      RECT 3.055 2.85 5.39 3.04 ;
      RECT 9.275 0.425 9.565 0.615 ;
      RECT 9.09 1.835 9.465 2.025 ;
      RECT 9.275 0.425 9.465 2.58 ;
      RECT 7.525 0.71 8.39 0.9 ;
      RECT 8.2 0.71 8.39 2.115 ;
      RECT 7.345 1.925 8.39 2.115 ;
      RECT 10.715 1.73 10.905 2.215 ;
      RECT 9.82 2.025 10.905 2.215 ;
      RECT 7.345 1.925 7.535 3.04 ;
      RECT 9.82 2.025 10.01 3.04 ;
      RECT 7.345 2.85 10.01 3.04 ;
  END
END XNOR3V2_7TV50

MACRO XOR2V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2V1_7TV50 0 0 ;
  SIZE 6.72 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.425 1.115 3 1.31 ;
        RECT 2.81 1.115 3 1.85 ;
        RECT 2.81 1.51 3.25 1.85 ;
        RECT 2.81 1.66 4.465 1.85 ;
        RECT 4.185 1.66 4.465 2 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.79 1.52 6.19 2 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.195 2.4 0.475 3.48 ;
        RECT 5.435 2.795 5.715 3.48 ;
        RECT 0 3.24 6.72 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.68 ;
        RECT 4.73 -0.12 5.01 0.565 ;
        RECT 0 -0.12 6.72 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.035 0.71 2.225 2.95 ;
        RECT 2.035 1.51 2.28 1.91 ;
        RECT 2.035 0.71 3.18 0.9 ;
        RECT 2.035 2.735 4.09 2.95 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 1.73 -0.24 3.505 1.545 ;
        RECT -0.12 -0.24 6.84 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 1.73 3.94 ;
        RECT 3.505 1.46 7.3 3.94 ;
        RECT -0.58 1.545 7.3 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 1.1 1.72 1.475 2 ;
      RECT 1.1 0.58 1.29 2.48 ;
      RECT 1.88 0.32 3.95 0.51 ;
      RECT 3.76 0.32 3.95 0.955 ;
      RECT 5.675 0.58 5.865 0.955 ;
      RECT 3.76 0.765 5.865 0.955 ;
      RECT 5.005 0.765 5.195 2.535 ;
      RECT 2.9 2.345 6.565 2.535 ;
  END
END XOR2V1_7TV50

MACRO XOR2V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2V2_7TV50 0 0 ;
  SIZE 8.16 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.36 1.52 6.605 1.995 ;
        RECT 6.36 1.8 7.22 1.995 ;
        RECT 5.99 1.805 7.22 1.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 1.52 1.32 2.005 ;
        RECT 0.54 1.81 1.77 2.005 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 2.405 0.435 3.48 ;
        RECT 1.865 2.79 2.145 3.48 ;
        RECT 5.515 2.79 5.795 3.48 ;
        RECT 7.315 2.4 7.595 3.48 ;
        RECT 0 3.24 8.16 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0.155 -0.12 0.435 0.735 ;
        RECT 1.955 -0.12 2.235 0.64 ;
        RECT 5.515 -0.12 5.795 0.66 ;
        RECT 7.315 -0.12 7.595 0.66 ;
        RECT 0 -0.12 8.16 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.99 0.71 4.18 1.395 ;
        RECT 3.94 0.71 4.22 0.91 ;
        RECT 3.99 1.205 5.11 1.395 ;
        RECT 4.92 1.205 5.11 2.595 ;
        RECT 3.565 2.4 5.11 2.595 ;
        RECT 4.92 1.995 5.16 2.32 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 2.475 -0.24 5.12 1.53 ;
        RECT -0.12 -0.24 8.28 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 2.475 3.94 ;
        RECT 5.12 1.46 8.74 3.94 ;
        RECT -0.58 1.53 8.74 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.92 0.71 3.2 1.42 ;
      RECT 2.76 1.215 2.955 2.64 ;
      RECT 3.405 0.955 3.595 2.08 ;
      RECT 3.405 1.89 4.68 2.08 ;
      RECT 2.435 0.32 5.135 0.51 ;
      RECT 4.945 0.32 5.135 0.66 ;
      RECT 1.1 0.595 1.29 1.03 ;
      RECT 1.1 0.84 2.625 1.03 ;
      RECT 2.435 0.32 2.625 1.035 ;
      RECT 2.335 0.84 2.535 2.55 ;
      RECT 1.06 2.36 2.535 2.55 ;
      RECT 1.06 2.36 1.25 2.79 ;
      RECT 2.345 0.84 2.535 3.035 ;
      RECT 4.415 2.795 4.695 3.035 ;
      RECT 2.345 2.845 4.695 3.035 ;
      RECT 6.46 0.595 6.65 1.195 ;
      RECT 5.45 1.005 6.65 1.195 ;
      RECT 5.34 1.61 5.64 1.8 ;
      RECT 5.45 1.005 5.64 2.43 ;
      RECT 5.45 2.24 6.68 2.43 ;
  END
END XOR2V2_7TV50

MACRO XOR3V1_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3V1_7TV50 0 0 ;
  SIZE 11.04 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.44 1.815 1.8 2.32 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.92 0.94 2.39 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.76 0.98 9.16 1.39 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.01 2.735 1.29 3.48 ;
        RECT 4.74 2.63 5.02 3.48 ;
        RECT 9.395 2.79 9.675 3.48 ;
        RECT 0 3.24 11.04 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.055 -0.12 1.335 0.615 ;
        RECT 4.895 -0.12 5.175 0.615 ;
        RECT 9.345 -0.12 9.625 0.615 ;
        RECT 0 -0.12 11.04 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.2 0.56 10.48 0.88 ;
        RECT 10.29 0.56 10.48 2.5 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 0.685 -0.24 8.625 1.565 ;
        RECT -0.12 -0.24 11.16 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 0.685 3.94 ;
        RECT 8.625 1.46 11.62 3.94 ;
        RECT -0.58 1.565 11.62 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 0.2 1.395 2.455 1.585 ;
      RECT 2.26 1.395 2.455 1.675 ;
      RECT 0.2 0.38 0.39 2.82 ;
      RECT 0.2 2.53 0.44 2.82 ;
      RECT 2.06 0.7 2.255 1.125 ;
      RECT 2.06 0.935 2.845 1.125 ;
      RECT 2.655 1.45 3.32 1.64 ;
      RECT 2.655 0.935 2.845 2.195 ;
      RECT 2.025 2.005 2.845 2.195 ;
      RECT 2.025 2.005 2.215 2.82 ;
      RECT 3.935 0.71 4.215 0.9 ;
      RECT 3.935 0.71 4.125 2.65 ;
      RECT 3.74 2.46 4.125 2.65 ;
      RECT 5.855 0.71 6.135 0.9 ;
      RECT 5.855 0.71 6.065 2.67 ;
      RECT 5.59 2.48 6.065 2.67 ;
      RECT 3.02 0.32 4.605 0.51 ;
      RECT 5.38 0.32 8.065 0.51 ;
      RECT 3.02 0.32 3.21 0.665 ;
      RECT 4.415 0.86 5.57 1.05 ;
      RECT 5.38 0.32 5.57 1.05 ;
      RECT 4.415 0.32 4.605 1.23 ;
      RECT 7.875 0.32 8.065 2.535 ;
      RECT 7.35 2.345 8.065 2.535 ;
      RECT 2.875 2.69 3.065 3.04 ;
      RECT 4.35 1.05 4.54 3.04 ;
      RECT 2.875 2.85 4.54 3.04 ;
      RECT 8.27 0.425 8.725 0.615 ;
      RECT 8.27 0.425 8.46 2.605 ;
      RECT 8.27 2.415 8.725 2.605 ;
      RECT 6.545 0.71 7.155 0.9 ;
      RECT 9.005 1.83 10.065 2.02 ;
      RECT 6.545 0.71 6.735 3.04 ;
      RECT 9.005 1.83 9.195 3.04 ;
      RECT 6.545 2.84 9.195 3.04 ;
  END
END XOR3V1_7TV50

MACRO XOR3V2_7TV50
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3V2_7TV50 0 0 ;
  SIZE 12.48 BY 3.36 ;
  SYMMETRY X Y ;
  SITE uhd50_CoreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.56 0.56 1.89 1.26 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.6 1.91 0.95 2.32 ;
        RECT 3.77 1.13 3.96 2.1 ;
        RECT 0.6 1.91 3.96 2.1 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.68 1.555 10.06 1.96 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.065 2.765 1.345 3.48 ;
        RECT 5.575 2.745 5.855 3.48 ;
        RECT 10.21 2.795 10.49 3.48 ;
        RECT 12.045 2.405 12.325 3.48 ;
        RECT 0 3.24 12.48 3.48 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.075 -0.12 1.36 0.73 ;
        RECT 5.605 -0.12 5.885 0.565 ;
        RECT 10.215 -0.12 10.495 0.615 ;
        RECT 12.045 -0.12 12.325 0.615 ;
        RECT 0 -0.12 12.48 0.12 ;
    END
  END VSS
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.155 0.53 11.4 0.88 ;
        RECT 11.205 0.53 11.4 2.65 ;
    END
  END Z
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER SN ;
        RECT 4.025 -0.24 9.115 1.53 ;
        RECT -0.12 -0.24 12.6 1.46 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER NW ;
        RECT -0.58 1.46 4.025 3.94 ;
        RECT 9.115 1.46 13.06 3.94 ;
        RECT -0.58 1.53 13.06 3.94 ;
    END
  END VNW
  OBS
    LAYER M1 ;
      RECT 2.135 1.295 2.85 1.485 ;
      RECT 2.135 1.295 2.325 1.685 ;
      RECT 0.21 1.495 2.325 1.685 ;
      RECT 0.21 0.54 0.4 2.58 ;
      RECT 2.09 0.54 2.28 1.095 ;
      RECT 3.38 0.74 4.445 0.93 ;
      RECT 2.09 0.905 3.57 1.095 ;
      RECT 4.255 0.74 4.445 2.545 ;
      RECT 1.96 2.355 4.445 2.545 ;
      RECT 1.96 2.355 2.15 2.82 ;
      RECT 4.645 0.71 4.925 0.9 ;
      RECT 4.695 0.71 4.885 2.65 ;
      RECT 4.695 2.46 4.975 2.65 ;
      RECT 6.48 0.71 6.845 0.9 ;
      RECT 6.48 0.71 6.67 2.82 ;
      RECT 7.785 1.1 8.11 1.41 ;
      RECT 6.87 1.205 8.11 1.41 ;
      RECT 6.87 1.205 7.06 2.125 ;
      RECT 2.99 0.32 5.365 0.51 ;
      RECT 6.085 0.32 8.89 0.51 ;
      RECT 2.99 0.32 3.18 0.705 ;
      RECT 5.175 1.335 6.275 1.525 ;
      RECT 6.085 0.32 6.275 2.105 ;
      RECT 8.7 0.32 8.89 2.565 ;
      RECT 8.15 2.375 8.89 2.565 ;
      RECT 2.765 2.745 3.045 3.04 ;
      RECT 5.175 0.32 5.365 3.04 ;
      RECT 2.765 2.85 5.365 3.04 ;
      RECT 9.275 0.425 9.565 0.615 ;
      RECT 9.09 1.055 9.465 1.255 ;
      RECT 9.275 0.425 9.465 2.61 ;
      RECT 7.585 0.71 8.5 0.9 ;
      RECT 8.31 0.71 8.5 1.87 ;
      RECT 7.345 1.68 8.5 1.87 ;
      RECT 10.715 1.73 10.905 2.49 ;
      RECT 9.82 2.3 10.905 2.49 ;
      RECT 7.345 1.68 7.535 3.04 ;
      RECT 9.82 2.3 10.01 3.04 ;
      RECT 7.345 2.85 10.01 3.04 ;
  END
END XOR3V2_7TV50

END LIBRARY
